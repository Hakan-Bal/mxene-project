H   8 A��@��\D�~��h��;M]�~F��)	��&��@��'3M]?[pQ)l�����1L��?)�Df��D@H            �         P   �������`���T������p���D����������̎����������l��������������f���񀄽�}�����P   P   ���䂄����z���;���<�������~�� ���y���V�����������~�������r���͇��]���ↄ�����P   P   �}������󂄽z���6�������S���ގ��*���#���ވ��S���V���Q�����������0�����������ↄ�P   P   񀄽5���B���8���߅������M~�����.�������������������U�������-���$����������]���P   P   f������鋄�[���ᄄ�S�������w������Y������`�����������0���v�������$���0���͇��P   P   ����H������m�����������̅��������������H�������G����|����������v���-�������r���P   P   ����񎄽���䅄�E���܊������������������l���_���^������ł������0���������������P   P   �������K������鉄��������4���1���6�������O����~��@�������|������U���Q���~���P   P   l���K���|���N��������������j���O�������ׄ����������~��^���G�����������V�������P   P   ����L���ኄ�����9���q���Ή��Q�������Ӎ������,������O���_�������`�������S�������P   P   ����B�������`���߄��)���K���Ո��č������D�������ׄ������l���H����������ވ��V���P   P   ̎��	�����������~��)���.������)���s�������Ӎ������6�����������Y�������#���y���P   P   ���匄�J���󅄽���ԋ��������l���)���č������O���1��������������.���*��� ���P   P   ����~���.�������l~������q|��Y���������Ո��Q���j���4�����������w������ގ���~��P   P   D���󎄽υ��ٍ��o���_������q|�����.���K���Ή�������������̅������M~��S������P   P   p���Ê������*����������_�������ԋ��)���)���q����������܊������S�����������<���P   P   ����胄�ފ��팄�,������o���l~������~��߄��9�������鉄�E�������ᄄ�߅��6���;���P   P   T������Ӂ��U���팄�*���ٍ������󅄽���`�������N������䅄�m���[���8���z���z���P   P   `�����������Ӂ��ފ������υ��.���J�����������ኄ�|���K���������鋄�B���󂄽���P   P   ����Ԁ����������胄�Ê��󎄽~���匄�	���B���L���K�������񎄽H������5�������䂄�P   P   �����������́��y����������|���3|��zq���z��u���v������|������򀄽����s������P   P   �������F|��}��F��x��p|���}�����w��/���{��z������{��n|���}��Gz���}��f~��P   P   s������@����|���~�������ey��&y���w��,|���z���x��z���x���{���~�� �W~���}��P   P   ���������|������7���}��ꁄ��|���z�����=����u���z�������|�������|����� �Gz��P   P   򀄽�����s��K������$|���|���{��<~���{��)�����L}��S���|��\|��Qx���|���~���}��P   P   ����j����z�����I���}���}���|���}�����t��~�����������|���x��\|�������{��n|��P   P   |��ly���|��}���z���|���{��~��Ex���{��}��V~��݀��]�������|��|���|���x���{��P   P   ����y��(t��|���x��\u��@z��X���m����{��y��-~��݅������]�������S�������z�����P   P   �v��z������|������{���{��w{��6x���v��D|���z��|��݅��݀������L}���z���x��z��P   P   u��Rr��8��}���v���y��M|���|��_u���s���z���y���z��-~��V~��~������u���z���{��P   P   �z��3~���y�� z��r|��a������F|���z�� z�������z��D|��y��}���t��)��=���,|��/��P   P   zq��lz�����Px��$���8���~�����~���{�� z���s���v���{���{�����{������w���w��P   P   3|���r��y}��fz��؀��{��[t���{��|��~���z��_u��6x��m���Ex���}��<~���z��&y����P   P   |���Sz��m{��|�����~��8���F����{����F|���|��w{��X���~���|���{���|��ey���}��P   P   ����ew��0����y��<���Lz��/x��8���[t��~������M|���{��@z���{���}���|��ꁄ��p|��P   P   ����Hw���u��*{���x������Lz��~��{��8���a����y���{��\u���|��}��$|���}������x��P   P   y�������w��W���z���x��<������؀��$���r|���v������x���z��I�������7���~��F��P   P   ́�������9z��W��*{���y��|��fz��Px�� z��}���|��|��}�����K�������|��}��P   P   ����}���w�����w���u��0���m{��y}������y��8�����(t���|���z���s���|��@���F|��P   P   ���������}���������Hw��ew��Sz���r��lz��3~��Rr��z��y��ly��j������������������P   P   y���p��Zr���v���t���w���t��p���v���~���v���{���z��q��v���v��;t��pq���r��p��P   P   p��Nr��nr���u���s���t���w���z��2y��4{��;x���s���|���v���{��;y���t��[t��u���v��P   P   �r���n��aq��w��s��!r��u��t���w��ax��1{���y��c~���u���u��Nv��jn���v���t��u��P   P   pq���t���t��/r���u��'u���w���t���y���s���u���t���v��ou��u��Zx��}v���w���v��[t��P   P   ;t��9o���y��lu���o���u��2t���q���z��2y���q��8v��&s���t���u��Fy��Gw��}v��jn���t��P   P   �v���r��ix��x��cp��\x���y���v��.w��Yw��ev���w��v��iu��zu���v��Fy��Zx��Nv��;y��P   P   v���t���z�� y��5u���w��u��-w��ty��Ru��Xw��{v���r��ao��]q��zu���u��u���u���{��P   P   q��cx���z��$v��2y���|���u��u��Vu���t���u���s��r��tr��ao��iu���t��ou���u���v��P   P   �z��7y��N|���u��Qx��Iz���y��Wz��Qz���|��$}���w���t��r���r��v��&s���v��c~���|��P   P   �{��u����t��*u��@z��cw���u���x���{��)}��ww��Ou���w���s��{v���w��8v���t���y���s��P   P   �v��Q~��$v��`s���v��zq��/r��is��bu���|���v��ww��$}���u��Xw��ev���q���u��1{��;x��P   P   �~���{���s���x��5{��u��
x��<z���v���w���|��)}���|���t��Ru��Yw��2y���s��ax��4{��P   P   �v������1s���w���t���o��+x��}q���u���v��bu���{��Qz��Vu��ty��.w���z���y���w��2y��P   P   p���z��Gx���t��D|��`l���~���y��}q��<z��is���x��Wz��u��-w���v���q���t��t���z��P   P   �t��9u��}��Sq���v��ex��mx���~��+x��
x��/r���u���y���u��u���y��2t���w��u���w��P   P   �w���x��{���|��t��fp��ex��`l���o��u��zq��cw��Iz���|���w��\x���u��'u��!r���t��P   P   �t��q���y���r���~��t���v��D|���t��5{���v��@z��Qx��2y��5u��cp���o���u��s���s��P   P   �v��l���z��y���r���|��Sq���t���w���x��`s��*u���u��$v�� y��x��lu��/r��w���u��P   P   Zr���u��~w���z���y��{��}��Gx��1s���s��$v���t��N|���z���z��ix���y���t��aq��nr��P   P   �p��*n���u��l��q���x��9u���z�������{��Q~��u���7y��cx���t���r��9o���t���n��Nr��P   P   Cm�� r��In���k���s���g���i���m��Uf���j���j���h��	k��ai���k���h���p��@m���m���p��P   P   �p���p���s���l���m���q���j��6j��ni���g��g���j��~g��ug���j���k���n���r���m���p��P   P   �m��Ds���m��dn��So���l���l���n���k���l���e��j��Zh���l��Lo��ul��o���j���k���m��P   P   @m��Gn���n��]k��&o��rm���l���l���l��=l���l��Ns��yn���h��Sp���g��o��n���j���r��P   P   �p��cp���p���o��q��m���n���q��5g��Xk��Tn���j��p��k���n���i��ti��o��o���n��P   P   �h���l��k��Kh���k���n���h���k��k��d��Ct��Xl��$k���l���o���n���i���g��ul���k��P   P   �k��an��jh��f���l���m��Rk���h���q���o���n��&m���l��}t���k���o���n��Sp��Lo���j��P   P   ai���o��1n���k��Hl���m��gl��In���g���i���i��0m���j���u��}t���l��k���h���l��ug��P   P   	k��[i��fc���g��ie��Wc��%e���h��Rg��i�� i��Dm���t���j���l��$k��p��yn��Zh��~g��P   P   �h��ch��3i��/n��$r��	q���o��k��lh���j��Jk��Pi��Dm��0m��&m��Xl���j��Ns��j���j��P   P   �j��g`��n���q���k���k���l��p��Am��8f���`��Jk�� i���i���n��Ct��Tn���l���e��g��P   P   �j���d��k���n��"e���i���j��j��k���j��8f���j��i���i���o��d��Xk��=l���l���g��P   P   Uf��Sh���m��|n��"k��v��~r���q���l��k��Am��lh��Rg���g���q��k��5g���l���k��ni��P   P   �m��0j��vj���n���e��^q���`���\���q��j��p��k���h��In���h���k���q���l���n��6j��P   P   �i���q���_���q���k��Tn���o���`��~r���j���l���o��%e��gl��Rk���h���n���l���l���j��P   P   �g��p��ej��_f���r���f��Tn��^q��v���i���k��	q��Wc���m���m���n��m��rm���l���q��P   P   �s���h���o��h��i���r���k���e��"k��"e���k��$r��ie��Hl���l���k��q��&o��So���m��P   P   �k��	p��!f��[j��h��_f���q���n��|n���n���q��/n���g���k��f��Kh���o��]k��dn���l��P   P   In��p���u��!f���o��ej���_��vj���m��k��n��3i��fc��1n��jh��k���p���n���m���s��P   P    r��bm��p��	p���h��p���q��0j��Sh���d��g`��ch��[i���o��an���l��cp��Gn��Ds���p��P   P   Z^��'a���f��Pa��c��9e���f��!k��9j��te��Sn���g���h���l���f��vf��`��Qe���b���b��P   P   �b���]���^���c��W`��$`��Fh���d��yh��}l���j��ym��6f��Qj��ld���d���b���a���b���_��P   P   �b���e��;e��d_���f��h��!e���f��Nb���h���e���e��ke��:h���e��d���i��:e��;d���b��P   P   Qe��|a��`��*g��ja���c���`��	c��ic��3f��^f���a���b��h��nd���c��_b���_��:e���a��P   P   `���d���Z���b���e���`��f���g��Ik��}f���e���c���b���f��ud���f��Go��_b���i���b��P   P   vf���j���h���i��%h���b��i���`��%e���h��l_���c���g��	f���c��^���f���c��d���d��P   P   �f��d���b��2i��$g��f`��Wf��Zh���`���f��wb���b��*f���_��d���c��ud��nd���e��ld��P   P   �l��b��na��n��!i���b���d���k���k��	h���g��Ve��ug��%^���_��	f���f��h��:h��Qj��P   P   �h��Kj���h���k��h��fi���k��j��6f��f���g��@b��pa��ug��*f���g���b���b��ke��6f��P   P   �g���c���i���e��U[��c��ie���d���e��j��j��Xh��@b��Ve���b���c���c���a���e��ym��P   P   Sn��m���e��[d���e��j���d��yc���e��l���n��j���g���g��wb��l_���e��^f���e���j��P   P   te��?k���k���^���b���f��c���b��g��g��l��j��f��	h���f���h��}f��3f���h��}l��P   P   9j��/c���g��*d���g��f���b��gf���b��g���e���e��6f���k���`��%e��Ik��ic��Nb��yh��P   P   !k���i���f���a��Ic��h��uj���p��gf���b��yc���d��j���k��Zh���`���g��	c���f���d��P   P   �f���d���h��i���d���c��Wb��uj���b��c���d��ie���k���d��Wf��i��f���`��!e��Fh��P   P   9e���_��mc���i��-`��lj���c��h��f���f��j��c��fi���b��f`���b���`���c��h��$`��P   P   c���k��;c��4p��`��-`���d��Ic���g���b���e��U[��h��!i��$g��%h���e��ja���f��W`��P   P   Pa���h��7e���h��4p���i��i���a��)d���^��[d���e���k��n��2i���i���b��*g��d_���c��P   P   �f���\��T^��7e��;c��mc���h���f���g���k���e���i���h��na���b���h���Z��`��;e���^��P   P   'a��Gh���\���h���k���_���d���i��/c��?k��m���c��Kj��b��d���j���d��|a���e���]��P   P   k��\���[��"b��fV��W`��]��oQ��Y��DX��+M��)X���W���T��\��E_��?Z���_��9[���^��P   P   �^��a��|^��'b���_��Y[��IZ��<Z��DW��X��7U��jS��?[��W��<Z���Y��`\���\��__���`��P   P   9[��+W���`���]��0Z���]��']��5\��e`��CV���]��]���\��TX��7\��O_���[���^���^��__��P   P   �_���c��s`���]��4_��5]��\��\��>\��U[���Z���]���]���\���V��]��hZ���[���^���\��P   P   ?Z��jY���b���Z���X��U^��y\��sX��Y��
Z��\��A^��8[���[��F]���\���Y��hZ���[��`\��P   P   E_��'W���Z���\��X��[��?_��H^���[��a��\��^��]���Z��c\���a���\��]��O_���Y��P   P   \���^���\��kW���X���c���Z���X��&[��X���[���^���]���\��ma��c\��F]���V��7\��<Z��P   P   �T��qX��t[���R��R��N[��|Y���N��,[��
Y���[���^���]��bY���\���Z���[���\��TX��W��P   P   �W��{W���^���\���\���_��*\���Y��Y���Y��J[��:_��LV���]���]��]��8[���]���\��?[��P   P   )X��\��UX���W���Y��g[���U��rZ���\���W��=S���[��:_���^���^��^��A^���]��]��jS��P   P   +M��[���Y��aZ���]��z]���Z��\��UZ��pV��9S��=S��J[���[���[��\��\���Z���]��7U��P   P   DX��TX���S���]���d���]��^��@c��]���T��pV���W���Y��
Y��X��a��
Z��U[��CV��X��P   P   Y���_���W���[��^^���O��<R���U��XZ��]��UZ���\��Y��,[��&[���[��Y��>\��e`��DW��P   P   oQ��/W���Z���[��Nd��ES��x^��Q^���U��@c��\��rZ���Y���N���X��H^��sX��\��5\��<Z��P   P   ]��LW��J_���R���\��mZ���X��x^��<R��^���Z���U��*\��|Y���Z��?_��y\��\��']��IZ��P   P   W`���^��$^���^���Z��-a��mZ��ES���O���]��z]��g[���_��N[���c��[��U^��5]���]��Y[��P   P   fV���Y���V���R���[���Z���\��Nd��^^���d���]���Y���\��R���X��X���X��4_��0Z���_��P   P   "b��qX��	`��$V���R���^���R���[���[���]��aZ���W���\���R��kW���\���Z���]���]��'b��P   P   �[��b���]��	`���V��$^��J_���Z���W���S���Y��UX���^��t[���\���Z���b��s`���`��|^��P   P   \���[��b��qX���Y���^��LW��/W���_��TX��[��\��{W��qX���^��'W��jY���c��+W��a��P   P   �G��&S���I��rQ���X���Q��+T���^��W���[���^��.Z���W��^Z��U��=Q���]���N��QS��dN��P   P   dN��qQ��(V���N���S��PY��O��SX��bZ��2T���\���Z��VY��XV��X��R���U���R���N��iV��P   P   QS��gS��dP��CR��cM���O��LS���N���U�� T��~V��]R��S���U���V���Q��Q���O���P���N��P   P   �N���P��0O��kL���V���S���V��QZ���T���V���T���R��{R��S��Y���U��X���Y���O���R��P   P   �]��S���S���V��Y��T���O��#V���O���R���T���R���X��T���S��nQ��M��X��Q���U��P   P   =Q��8Q��Q��aO���S��?R���L���V���T���Q���W��bQ���P���R��YQ��jU��nQ���U���Q��R��P   P   U���P��'\���[��~W��RU���V���T���Y���U���R��Q���P��(X���S��YQ���S��Y���V��X��P   P   ^Z���X��tV��!U��
]���R��CW���]��oV��bU��FS���S��gS��:[��(X���R��T��S���U��XV��P   P   �W���V���Q���O��(T���P��IN���W���X���W��$S��T���U��gS���P���P���X��{R��S��VY��P   P   .Z��V���T���W���^��ZV��@Y��<V���R��X��M^���R��T���S��Q��bQ���R���R��]R���Z��P   P   �^���T��X��rT���M��kL��mR��1V��3W��X���\��M^��$S��FS���R���W���T���T��~V���\��P   P   �[��KX��%W��GW��N��ZS���T���O���O��\��X��X���W��bU���U���Q���R���V�� T��2T��P   P   W���R��fV��>R���M��`���`��3Z���S���O��3W���R���X��oV���Y���T���O���T���U��bZ��P   P   �^���T��V���Y���N��aZ��XR��9K��3Z���O��1V��<V���W���]���T���V��#V��QZ���N��SX��P   P   +T���W��-Q���U���Q��_T���]��XR���`���T��mR��@Y��IN��CW���V���L���O���V��LS��O��P   P   �Q��}T��RT��6O���Y��K��_T��aZ��`��ZS��kL��ZV���P���R��RU��?R��T���S���O��PY��P   P   �X���P���Z���U��b[���Y���Q���N���M��N���M���^��(T��
]��~W���S��Y���V��cM���S��P   P   rQ��R���R���\���U��6O���U���Y��>R��GW��rT���W���O��!U���[��aO���V��kL��CR���N��P   P   �I���T���P���R���Z��RT��-Q��V��fV��%W��X���T���Q��tV��'\��Q���S��0O��dP��(V��P   P   &S��tT���T��R���P��}T���W���T���R��KX���T��V���V���X���P��8Q��S���P��gS��qQ��P   P   SL���P���O��6K��cI���H���F��$D��+H��?C��G���C���F��DF���I��QI��H��J���P���P��P   P   �P��YJ���J��\Q��CH��)I���T��I���E��LH��GC���E���D��I��I���R��UH���I���N���F��P   P   �P���T���L��MO��S���L���I���L��dC���M��5K��sJ��M��vJ��}D��WG���M���L���V���N��P   P   J��`G���L���L��YG��/O��}G���H��{L��J��FM���H��M��kK��K���K���H���G���L���I��P   P   H���O��-J��)O��H��zH��;M���I��vP���M���H��ZK���K��
M��eI���N��R���H���M��UH��P   P   QI��VN��fM��HJ��M���M��kR���J��I���L���J��'P��hN��L��|O���I���N���K��WG���R��P   P   �I���G��E���B��,H���A��<I��/H��tC���L���J���M���L��tE���H��|O��eI��K��}D��I��P   P   DF��JH���L���I��AM��cK���G��4J���C��UL��N��@L���J��1G��tE��L��
M��kK��vJ��I��P   P   �F��FJ��iI���I��yF��=H�� P��*H��3F���F��]K���J��sM���J���L��hN���K��M��M���D��P   P   �C���H��(L��,K��qI��kD���N��QH��_H���F���E��SH���J��@L���M��'P��ZK���H��sJ���E��P   P   G��E��AE��"L���O���O���P���G���G���G���A���E��]K��N���J���J���H��FM��5K��GC��P   P   ?C���G���L��NK���H��.H���F��F��mM���I���G���F���F��UL���L���L���M��J���M��LH��P   P   +H��LE��FI���L���K��[I��
G��H���R��mM���G��_H��3F���C��tC��I��vP��{L��dC���E��P   P   $D��L��YI��fF���H��jJ���B���I��H��F���G��QH��*H��4J��/H���J���I���H���L��I��P   P   �F���H���M��1P��N��:M��$B���B��
G���F���P���N�� P���G��<I��kR��;M��}G���I���T��P   P   �H��[G���I��WH��G���K��:M��jJ��[I��.H���O��kD��=H��cK���A���M��zH��/O���L��)I��P   P   cI���N���G���L���D��G��N���H���K���H���O��qI��yF��AM��,H��M��H��YG��S��CH��P   P   6K���R���G���B���L��WH��1P��fF���L��NK��"L��,K���I���I���B��HJ��)O���L��MO��\Q��P   P   �O���G���K���G���G���I���M��YI��FI���L��AE��(L��iI���L��E��fM��-J���L���L���J��P   P   �P��*Q���G���R���N��[G���H��L��LE���G��E���H��FJ��JH���G��VN���O��`G���T��YJ��P   P   K��J;��E���C���>���D��3G��DA���I��I��3G���J��<H���B��iD���F��>��{I��|?���?��P   P   �?��L@��=��x?��zC��qA���@��{E��H���I���E���F��F���K��DC��=?���B���B���A���9��P   P   |?��]8��<A���=��T<���F���A��SF���H��D���A���I���D��|D���H���G���E��C���8���A��P   P   {I���A���C���I���A���A���D���@���B��ZC��=B���E���B���B��VA���C��KB���@��C���B��P   P   >��G@���B��w:��8?��HB���A���C���@���A��C���D��,>��A���D��'@���?��KB���E���B��P   P   �F��qB��yF���G���C���F���A��D���D���B��<@��BA���B���C���B��B��'@���C���G��=?��P   P   iD���J��A���C���F��J��2A���E���G��+B��0C���C���C���I���F���B���D��VA���H��DC��P   P   �B���C���D��E���<��/E��!F���B��*M���D���>��4C��D��zG���I���C��A���B��|D���K��P   P   <H��;C���D��aH���M���D���E��y@��G��G���D���B��A��D���C���B��,>���B���D��F��P   P   �J���I���C��<���<���A���;���A���L���J��KE��K���B��4C���C��BA���D���E���I���F��P   P   3G��K���C���B��#D���D��UE��GB��H��+G���G��KE���D���>��0C��<@��C��=B���A���E��P   P   I��E���@��0?��I��E��BG���E��nD��m:��+G���J��G���D��+B���B���A��ZC��D���I��P   P   �I���L��F���D���G��{<���?���?��(B��nD��H���L��G��*M���G���D���@���B���H��H��P   P   DA��hD��B���>��uG��"B��Q���S���?���E��GB���A��y@���B���E��D���C���@��SF��{E��P   P   3G�� F��@���?��DC��/A���C��Q���?��BG��UE���;���E��!F��2A���A���A���D���A���@��P   P   �D��TJ���C���G��;C���F��/A��"B��{<��E���D���A���D��/E��J���F��HB���A���F��qA��P   P   �>��5C���@���D���D��;C��DC��uG���G��I��#D���<���M���<���F���C��8?���A��T<��zC��P   P   �C���>���G��]D���D���G���?���>���D��0?���B��<��aH��E���C���G��w:���I���=��x?��P   P   E���A��E���G���@���C��@��B��F���@���C���C���D���D��A��yF���B���C��<A��=��P   P   J;���9���A���>��5C��TJ�� F��hD���L��E��K���I��;C���C���J��qB��G@���A��]8��L@��P   P   �3���<��;���8���A��B9���7��?��/��76���6���3��25���=��2:���:��@>���6��F<���:��P   P   �:���A��eD��9��?��|>���1��a8���7���5���;��`8���7���1��59���1��f>��+>���;��-I��P   P   F<���;�� ;���;��::���6���;���7���8��e6��A7���5���5���7���7��q:���6��]=���5���;��P   P   �6��f?���<���6���A��8��I<��g?���8��(<���9���<���8���=���;���8��>���:��]=��+>��P   P   @>���6��w<���8��A?���>���8��=���8���=���>��<��?��E>���>��=���:��>���6��f>��P   P   �:��97���3��6���6��6��$5���8���:���;��7>��:��M9���<���6���=��=���8��q:���1��P   P   2:���4��#>��>C�� 9���6��T9���8���7��.;���>��':��7���6���5���6���>���;���7��59��P   P   �=���8��$1���7���5���3���:��<��s4�� 6��Z=�� =��R:���8���6���<��E>���=���7���1��P   P   25���8��m<���4���7��P;��7���:��$5��05��`9���:���;��R:��7��M9��?���8���5���7��P   P   �3���.���8��#A���=���@��=��z<���/��W1��8��6���:�� =��':��:��<���<���5��`8��P   P   �6���5��@��z:���6��1���3���<���:�� 5��^<��8��`9��Z=���>��7>���>���9��A7���;��P   P   76��3���:��8��7���:��;���8���7��>�� 5��W1��05�� 6��.;���;���=��(<��e6���5��P   P   /���2��:���6���5��=��L9��-=��h5���7���:���/��$5��s4���7���:���8���8���8���7��P   P   ?��&7���=���?���7���8��r.���'��-=���8���<��z<���:��<���8���8��=��g?���7��a8��P   P   �7���9���7���;��97���8���;��r.��L9��;���3��=��7���:��T9��$5���8��I<���;���1��P   P   B9���4��j6��3<��l:��m7���8���8��=���:��1���@��P;���3���6��6���>��8���6��|>��P   P   �A��j7��:��o6��;6��l:��97���7���5��7���6���=���7���5�� 9���6��A?���A��::��?��P   P   �8��N5���7���@��o6��3<���;���?���6��8��z:��#A���4���7��>C��6���8���6���;��9��P   P   ;���?���6���7��:��j6���7���=��:���:��@���8��m<��$1��#>���3��w<���<�� ;��eD��P   P   �<��1>���?��N5��j7���4���9��&7���2��3���5���.���8���8���4��97���6��f?���;���A��P   P   8*���2��g)���/���,���3��^2���3��?7��x:��"4��`8��z;���0���4���0��A0���*��6,�� 0��P   P    0���-���)���2���+���,���=���3���3��>7���1��4��:��S/���7���;��-��5/���/���*��P   P   6,��b5��?,��p3���9���.���3��_5��"1���9��R8���3��8���8���4��Q4���2��/���9���/��P   P   �*��;.���-���*���(��q2���.��b.��"3��2���3�� 3��#4���1���2��A/���0���/��/��5/��P   P   A0���:��3��.<���/���-��I6���-��	5��1��v,���-��B0���/���)��@2���4���0���2��-��P   P   �0���7��t.��p/���7��1���9��4��2���0��/���7�� 5���4��\7���1��@2��A/��Q4���;��P   P   �4���0��C4��+���1��U2��	8��5��V4���2���-���2��R:��L4��*9��\7���)���2���4���7��P   P   �0��v1���;���4���8���:���/��s.��>0��~7���3��L/���3��7��L4���4���/���1���8��S/��P   P   z;��&6��
3��K0���'��2���.���6���<��|;���6���2���3���3��R:�� 5��B0��#4��8��:��P   P   `8���7��a-��x1���5��T0��1��f3���6��)8���3���0���2��L/���2���7���-�� 3���3��4��P   P   "4��k3���2��(.��h4���6��i4���1��,���5��95���3���6���3���-��/��v,���3��R8���1��P   P   x:���:���3���6���/��^0��R/���1��X2���:���5��)8��|;��~7���2���0��1��2���9��>7��P   P   ?7���6���.���2��5��7���7���5���4��X2��,���6���<��>0��V4��2��	5��"3��"1���3��P   P   �3���7��s0���0���2��;2��S7��7���5���1���1��f3���6��s.��5��4���-��b.��_5���3��P   P   ^2���0���3���-��o2��S4���5��S7���7��R/��i4��1���.���/��	8���9��I6���.���3���=��P   P   �3���2���7��y2��
2��75��S4��;2��7��^0���6��T0��2���:��U2��1���-��q2���.���,��P   P   �,���5��6��+2��1��
2��o2���2��5���/��h4���5���'���8���1���7���/���(���9���+��P   P   �/��(:��0���+��+2��y2���-���0���2���6��(.��x1��K0���4��+��p/��.<���*��p3���2��P   P   g)��$.���3��0��6���7���3��s0���.���3���2��a-��
3���;��C4��t.��3���-��?,���)��P   P   �2���0��$.��(:���5���2���0���7���6���:��k3���7��&6��v1���0���7���:��;.��b5���-��P   P   N2���+���1���1���%��)���'��M$��e(��s!���&���#���"��n%���&��f(��%���3��u/���-��P   P   �-��`&���&���)���+���*���#���%���(��$��u&��n)������,���#��_%���*���+���,��*#��P   P   u/��L*��|1���,��y"���0���&���%��>+��a$��r$���,���#��~$��b,��"���-��u(��c$���,��P   P   �3���%���'��C5���(���*��v-��[(���+��`*���*���(��,��B)���,���+���)��.��u(���+��P   P   %���&��z!��e!���)��[,��9)��?,���-��m*��/��C/��/+��?.��t/��+��u+���)���-���*��P   P   f(���%���/���/��%���(��# ���#���*��
,��R.���(���(���%��
*���,��+���+��"��_%��P   P   �&��*������'��A$��L'��M(���'��-���(��m1��<*���"���)��^%��
*��t/���,��b,���#��P   P   n%���'���(��)���'���&��c)��5%��G+���%���&��r-���(��.'���)���%��?.��B)��~$���,��P   P   �"���%��A$��Y,��r1��`)��J(���$���"��� ��e$��3*���,���(���"���(��/+��,���#�����P   P   �#��	+��
.��8$��%��e$���%��+��*���"��(��q0��3*��r-��<*���(��C/���(���,��n)��P   P   �&��$&���#��a-��M(��|*��@,��]*��C&���'���$��(��e$���&��m1��R.��/���*��r$��u&��P   P   s!���(��#��+'���*�� &�� &��[)��f(���$���'���"��� ���%���(��
,��m*��`*��a$��$��P   P   e(���$��E)��$)��(������"��B���(��f(��C&��*���"��G+��-���*���-���+��>+���(��P   P   M$���&���(��b*���)���"���'���+��B��[)��]*��+���$��5%���'���#��?,��[(���%���%��P   P   �'���&���(��*��3*���$��O#���'���"�� &��@,���%��J(��c)��M(��# ��9)��v-���&���#��P   P   )���*��P%���%��<)��%���$���"����� &��|*��e$��`)���&��L'���(��[,���*���0���*��P   P   �%���#��p%��]*���-��<)��3*���)��(���*��M(��%��r1���'��A$��%���)���(��y"���+��P   P   �1��{'��.*��e*��]*���%��*��b*��$)��+'��a-��8$��Y,��)���'���/��e!��C5���,���)��P   P   �1��&��m&��.*��p%��P%���(���(��E)��#���#��
.��A$���(������/��z!���'��|1���&��P   P   �+���)��&��{'���#���*���&���&���$���(��$&��	+���%���'��*���%���&���%��L*��`&��P   P   X����������)&���"��7%��a%���%���#���$��%������)���!���%��� �����������P   P   ���X���%�����!���#�����'��E#��b)���(��#'���)��]*���#������$�����r���"��P   P   ��� ��������������!���&�� $���!���&��� ��b&��Z"������&�����^"��
��r��P   P   ���b%��c(��8���#�����
��%��(��z!���#���������$�����k%���!��j��^"�����P   P   � ����6&����V ���&�����9$������q"��"���$���!��$�����q���!������$��P   P   �%��\"��� ��^!��	"��Z$��"���'��t ������ ��p��9'���%�����7 �����k%���&�����P   P   �!���$���"���'��m$��5#��� ��D$��\��!��� ���"��'��[)���&�����$���������#��P   P   �)���&���������������&���)��%��?%��N'��� ���'��c&��[)���%���!���$��Z"��]*��P   P   ���!���!��< ��8"���!��E%�� ���#���'��&��!��x���'��'��9'���$�����b&���)��P   P   %��I��X$���$�����3"��L#��� �� !��}&��P&�����!��� ���"��p��"������ ��#'��P   P   �$���&��_ ��� �����|��������o&��#���&��P&��&��N'��� ��� ��q"���#���&���(��P   P   �#��� ���'������ ��~'��@&������ ���!��#��}&���'��?%��!�������z!���!��b)��P   P   �%��!��7&��i ��� ���&���%���'��$��� ��o&�� !���#��%��\��t ����(�� $��E#��P   P   a%��� ���"��{��z��-+��n������'��������� �� ���)��D$���'��9$��%���&��'��P   P   7%��S%��j$��y#��Y ��%&��f%��n���%��@&�����L#��E%���&��� ��"�����
���!�����P   P   �"��	"��[ ��=��������%&��-+���&��~'��|��3"���!�����5#��Z$���&��������#��P   P   )&��#��������F�����Y ��z��� ��� ��������8"�����m$��	"��V ���#�����!��P   P   ��(��P#��#�����=��y#��{��i ������ ���$��< ������'��^!����8��������P   P   ����#��,#��P#�����[ ��j$���"��7&���'��_ ��X$���!������"��� ��6&��c(������%��P   P   ������#��(��#��	"��S%��� ��!��� ���&��I��!���&���$��\"����b%�� ��X��P   P   ���������}����������A������������g�������&��������l�����P   P   ���u"�����'�����z��Q��I�����Z��i����������0�����������G�����P   P   l��y��>����&�������� ������F��M��'�����x��������V��� ��G��P   P   ������������������������������������6��W�����b�������V�����P   P   ������t���!��n��C��������h��"����C��������������a�����������P   P   &��}������	��(��L�����������0!�����&��������d��y�����b��������P   P   �����������������A����E�����x��������������d��������x��0��P   P   ���������J��m�����6�����u�����B�����!�������������W��������P   P   g��L��R����D����]��v�����������c��4��!�����������6��'����P   P   ���S�����,�����x�����/�����u��%��|��c��������&��C�����M�����P   P   ��B�����������m��~��"�����������%�����B��x����������F��i��P   P   ����p��<��X��-��!�����M��!�����u�����������0!��"�������Z��P   P   ���H����#��?�������=����M�����������u��E�����h����������P   P   A��������Y��-�����������=�����"��/��v���������������� ��I��P   P   �����������������������!��~�����]��6��A��������������Q��P   P   ���H�����������������������-��m��x����������L��C��������z��P   P   ���H��������4�������-��?��X��������D��m�����(��n�����&�����P   P   }�����i��������������Y��#��<�����,����J������	���!�������'��P   P   ��������i����������������p��������R�����������t�����>�����P   P   ���]��������H��H��������H����B��S��L��������}��������y��u"��P   P   �����$��.��w��M��������T�����������w�����h��n������������
��P   P   �
�������h���������������������z��������������������L
��P��P   P   ���������~��g ���������������E��9��E��y��������x��2��E��L
��P   P   ���\��6�����
���������?��Q��9��������@�����i��U��s��2�����P   P   ���������������������:������
�����%�����D�������D��U��x�����P   P   n���
���������
���������	�����
��b�����I��^��q��������i��������P   P   h�����%����D
��J��������[�������������������q�������������P   P   ��������A��!��������������y��$�����C��" �����^��D��@��y�����P   P   w�����|��������o��x�����������������p��C�����I��������E�����P   P   ���J��Y����������z�����i��O��2�����������������%�����9��z��P   P   ������������l����K��*��b�������2�����$����b�����9��E����P   P   ���!��T������������������������O�����y�����
���
��Q��������P   P   T�����m��a�����D��������3����b��i��������[��������?��������P   P   ���������m��������������������*���������������	��:���������P   P   ������0�����������������������K��z��x����������������������P   P   M�����������;�����������D���������o�����J���������������P   P   w��f�����������;��������������l��������!��D
���
������
��g �����P   P   .�����a��)�����������m��a��������������A������������~��h��P   P   $�����~��a��������0�����m��T�����Y��|�����%��������6�������P   P   ��T��������f��������������!�����J�����������
�����\��������P   P   1�����	��X ������������>��U	���������u������������������A����u
��P   P   u
��� �����.����������������q��������������������H��		���
�����P   P   ��G������
��@
��;�������C�����������J���������W
�����<���
��P   P   A����a
��k����� �� ��
��P�����X��N��F	������������	��������		��P   P   ���� �����������a�������2�������������D��_��@������	��W
��H��P   P   ��������q	��������������4��v��L��+��f��
��E��e��@�����������P   P   ����������)��q�����u�����������������������O��E��_����������P   P   ���7������������/��� �����r��<��
����������
��D�����������P   P   �������T
���
��������� ��^��8
��J��R��m
��������f�����F	��J����P   P   u�����U��c�����	�����r�����������b��R��
�����+�����N��������P   P   ����������� ��� �����i���+��Q�����������J��<�����L�����X��������P   P   ���0
���
������c����_������6�����������8
��r�����v����������q��P   P   U	�����5��;��6�����e�����m ��6��Q�����^��������4��2��P��C�����P   P   >�����b��5 ��� ��������������������+��r��� ��� ����������
�������P   P   ����W������������v��������e��_��i���������/��u�������� �������P   P   ����	�����L�����_��v�������������	��������������a�� ��;�����P   P   ������t��9�� 	���������� ��6��c��� ������
����q����������@
�����P   P   X �����3��5��9��L�����5 ��;������� ��c��T
����)��q	������k���
��.��P   P   	��������3��t��������b��5���
�����U����������������a
��������P   P   ���b������������	��W��������0
����������7�������� ����G��� ��P   P   ����"�=���g���������������	�����������%��|�����g������s����󃽞���P   P   ����4�������􃽿�������� ��6������������������X���X����x���Y���I���3��P   P   ������X���|���� ��R��������� �����9��������������~����������I���P   P   s�����������������������* ��:���������$��:
��W��c��[�������������Y���P   P   ���� ��>������G���������������������f���������T���m��c������������x���P   P   g����������q�����������������������������V��f
����0��c��[���~����P   P   �������k ���������S���k�����( ���������	��<����������m��c������X��P   P   |��`������ ����������d��+������D�����R����
�� �����f
��T���W����X���P   P   %������ �������������������������� ������
���
��<��V����:
��������P   P   ���B��I������G����������.���G ����2��1�����R���	���������$��������P   P   ���� �����,�������������������������2�� ������������f������9�����P   P   ����������f��� ������9���Q�� ����������������D��������������������P   P   	���������� ��G ���������<������� ������G ���������( ����������:���� ������P   P   ���Q��,������e��F������� ��<���Q����.������+������������* ����6��P   P   ���. ����������������� ���������9��������������d��k��������������� ��P   P   ������� �����������������F��������������������������S���������������R�������P   P   ������Z���~������������e��G ��� �����G����򃽔���������G������� ������P   P   g���W ��<���� ��~��������������� ��f��,���������� ������q���������|�����P   P   =�����������<���Z��� ������,��������������I���� �����k ������>������X������P   P   "�K�������W ���������. ��Q��������� ��B�����`���������� ����������4���P   P   �샽����C�����󃽸󃽒򃽀������������0􃽅��������_�������B�P   P   B񃽱���P����􃽰��������������������[���z��������������3���z���'�������P   P   ����5���k���O���9���y3����샽���������}�����������V����&�n���n􃽞�P   P   _���0탽?샽���������󃽃���������������Q���q���[���������������H�������n���'���P   P   ��/���H󃽜���������������x������������������H���&�z���P   P   ��4ꃽ��������m�������2[�������A�������􃽼���c���q�����������3���P   P   �������������������������@�������� ������c ������c����������V������P   P   �p��􃽏����􃽕������������������!������c ���������������������P   P   0��h�����������#����􃽾􃽈񃽶�������������!�������������[�����������P   P   ��������c��������������������g���������� �����x��q���}���z���P   P   ����������탽8��������� ���������������A�����Q�����[���P   P   �Z�������!��zcj򃽥샽M�������򃽶�������@����������������������P   P   ���������M7ꃽ�������샽�����󃽈��������[�����������������P   P   ��h��󃽵�탽L�都�僽�j򃽏�򃽾�����2��������샽��P   P   �򃽃�B�r���t����都��c8���������������������3�������P   P   ���񃽠���$�����2샽��L��z탽��#�������m���H���y����P   P   󃽫냽{���3������􃽴�탽7ꃽ�����������������9�������P   P   �����탽2���s���3�$���r�M!��c������������������������O�����P   P   C���2���{�������B��������������h����􃽗�������?샽k���P���P   P   ����������탽�냽�񃽃�h󃽾�Z�����������p󃽬���4ꃽ/0탽5�������P   P   �能�能"⃽c能�⃽��탽����������"탽H񃽿���T���냽�K都'烽�惽n惽P   P   n惽3ჽ2⃽/냽�都�E������������탽����􃽳������񃽒z샽�䃽⃽P   P   �惽yヽ'ヽ�能�惽U�탽����1�%�������������M����1�������烽�탽�䃽P   P   '烽�都�都f샽�惽*���D能yꃽY���샽����d�����������������탽�都�烽z샽P   P   K都都��烽�能�냽�,냽������������o���� ���������샽�탽����P   P   ��都�烽T䃽&샽_����탽'�����������|������ ����������󃽗���1�����P   P   냽S����ꃽmჽ�R�7�����Y􃽚냽���^����������.�����������������P   P   T����샽�탽䃽"ꃽ�能�탽�����t���� ��H���e������ ��� ������M��P   P   ����}���n烽能�烽�ヽi냽?����-�������y�������H���������o������������P   P   H񃽙񃽶�h샽�烽v惽S탽탽����L�h����y���� ��^���|�������d�����������P   P   "탽�탽�ꃽ�샽�ꃽ�냽hy탽�냽~ꃽh����t����������������������탽P   P   ����Y���1f냽�냽�샽M都O都`����都~L�-�����냽�����샽%�����P   P   �����탽�냽Kj����ꃽF샽�都`����냽�������Y�����Y���1���P   P   �����탽�냽r탽?탽;都@��都O都y탽탽?�������'���,냽zꃽ��������P   P   �탽�샽6샽��냽Kꃽ(ꃽ;都F샽M都hS탽i냽�탽7����탽�D能�탽E�P   P   �*�-都]ヽ�都HꃽKꃽ?탽�ꃽ�샽�냽v惽�ヽ�能R�_����냽*���U�P   P   �⃽�G샽�都烽�都�냽r탽j����냽�ꃽ�烽�烽"ꃽ�&샽�能�惽�惽�都P   P   c能?냽j僽;����都]ヽ��냽Kf냽�샽h샽能䃽mჽT䃽�烽f샽�能/냽P   P   "⃽�都�j僽G샽-都6샽�탽�냽1�ꃽ��n烽�탽�ꃽ�烽��都'ヽ2⃽P   P   �能ヽ�都?냽�*􃽪샽���탽Y����탽��}����샽S����都都�都yヽ3ჽP   P   �ۃ�
݃��ރ��܃��䃽�܃�7⃽:烽�⃽�샽��8ރ�4탽����A܃��僽�܃�݃�����P   P   �����܃�I烽Sჽ����ჽD݃�	냽hჽx能
ꃽ탽烽�ჽTꃽ����4߃��ۃ��ჽ�ヽP   P   ݃��܃�iჽ߃�S܃�Q能`ヽ�能K샽�탽�K惽p��能�䃽能W僽�ヽ�ჽP   P   �܃�=݃�߃��ۃ�ރ��烽�샽�샽�샽d�������I���������5탽.能�W僽�ۃ�P   P   �僽⃽�ڃ�B����僽h䃽MჽT`ꃽ���#�能�,能탽����v.能能4߃�P   P   A܃��⃽.ك�m܃�Bჽ ݃�����>都e냽��������F�����%���!�����������5탽�䃽����P   P   ����V؃�ヽ�僽}⃽�ԃ��ჽ�都G惽1�����z��������]���!���탽�����能TꃽP   P   4탽⃽�ۃ�惽�䃽)ރ��⃽�烽ヽ��j�_都I���>烽�%���,能������ჽP   P   8ރ�⃽�߃����ჽB߃�C僽_߃��ჽO僽���I������������I�p烽P   P   �D݃��߃��߃��݃��܃�m߃��݃�*ჽ�샽.都�탽�_都z���F򃽣能��K惽탽P   P   �{僽�����ރ��܃�mރ�s݃��ۃ��ჽ�ヽ��.都�j􃽣�����#���
ꃽP   P   �샽�ヽv߃�z܃��ۃ�=ك��ڃ��փ��ރ��܃��ヽ�샽O僽��1����������d����탽x能P   P   �⃽⃽S����܃��ڃ��Ӄ��Ӄ�Dك�ڃ��ރ��ჽ*ჽ�ჽヽG惽e냽`ꃽ�샽K샽hჽP   P   :烽Bރ�5߃��݃�*ك�؃�.܃�x݃�Dك��փ��ۃ��݃�_߃��烽�都>都T�샽�能	냽P   P   7⃽ヽ%䃽yჽ-܃�v׃��ڃ�.܃��Ӄ��ڃ�s݃�m߃�C僽�⃽�ჽ����Mჽ�샽`ヽD݃�P   P   �܃��؃�O݃��ރ��݃�rჽv׃�؃��Ӄ�=ك�mރ��܃�B߃�)ރ��ԃ� ݃�h䃽�烽Q能�ჽP   P   �䃽�䃽J����能�܃��݃�-܃�*ك��ڃ��ۃ��܃��݃�ჽ�䃽}⃽Bჽ�僽ރ�S܃����P   P   �܃��⃽�ك��烽�能�ރ�yჽ�݃��܃�z܃��ރ��߃����惽�僽m܃�B����ۃ�߃�SჽP   P   �ރ��ރ��׃��ك�J���O݃�%䃽5߃�S���v߃������߃��߃��ۃ�ヽ.ك��ڃ�߃�iჽI烽P   P   
݃�ރ��ރ��⃽�䃽�؃�ヽBރ�⃽�ヽ{僽D݃�⃽⃽V؃��⃽⃽=݃��܃��܃�P   P   σ�̓�Ѓ�҃�Ճ��ރ�����ރ��ჽ*ރ��׃��ރ��⃽�ك�)ჽ߃��ԃ�.Ճ�/у��˃�P   P   �˃�tσ��Ƀ�у��׃��ރ�-⃽ჽl냽�惽N�都e냽�都.���S⃽�݃��Ճ��Ӄ�Mȃ�P   P   /у�iӃ�9Ѓ��Ӄ�4ڃ��҃�&ރ��ރ�惽A냽D僽�탽e⃽�僽t���ۃ��؃��Ӄ��Ӄ�P   P   .Ճ�TЃ�Ѓ��σ��ۃ��Ճ��ك�mꃽ�݃� 탽'냽+�����?탽�能c僽�惽�փ��؃��Ճ�P   P   �ԃ�fЃ�(Ӄ�6҃��у��܃�6ك�D能�烽�냽	����,��������󃽻䃽J냽�惽ۃ��݃�P   P   ߃��҃��փ��ك��ԃ��܃��ヽ"⃽�⃽2都�탽���������\񃽻䃽c僽t���S⃽P   P   )ჽ�؃��ԃ��у�rу��ރ��߃�����䃽{샽I��������-����������󃽟能�僽.���P   P   �ك�I܃��׃�Ã�Uȃ�,ك�`܃� ۃ�8都n탽D탽E�����/���-���񃽉���?탽�都P   P   �⃽�܃�]ރ��Ճ��Ӄ��׃��׃��ڃ��烽3烽�ヽ����x����􃽢����,�����e⃽e냽P   P   �ރ�ჽ�׃��Ӄ�փ��փ��Ӄ�ڃ�R���'܃�7ꃽ�����E��������������+����탽�都P   P   �׃�ۃ��⃽�Ӄ��҃�G΃�F҃��փ��⃽�؃��݃�7ꃽ�ヽD탽I�탽	�'냽D僽NP   P   *ރ�Cك�6ރ��׃�O؃�׃��؃�ڃ�ԃ�߃��؃�'܃�3烽n탽{샽2都�냽 탽A냽�惽P   P   �ჽ�䃽b���2փ�yՃ�`ۃ�'փ��׃�]փ�ԃ��⃽R����烽8都䃽�⃽�烽�݃�惽l냽P   P   ރ��ڃ�tك��؃��ك��Ճ�-҃�WɃ��׃�ڃ��փ�ڃ��ڃ� ۃ�����"⃽D能mꃽ�ރ�ჽP   P   �����ރ�N؃��Ѓ�=҃��׃��҃�-҃�'փ��؃�F҃��Ӄ��׃�`܃��߃��ヽ6ك��ك�&ރ�-⃽P   P   �ރ�3ڃ�_ڃ��ڃ�GՃ�LӃ��׃��Ճ�`ۃ�׃�G΃��փ��׃�,ك��ރ��܃��܃��Ճ��҃��ރ�P   P   Ճ�#у�[у�;ȃ�׃�GՃ�=҃��ك�yՃ�O؃��҃�փ��Ӄ�Uȃ�rу��ԃ��у��ۃ�4ڃ��׃�P   P   ҃��Ѓ��܃��҃�;ȃ��ڃ��Ѓ��؃�2փ��׃��Ӄ��Ӄ��Ճ�Ã��у��ك�6҃��σ��Ӄ�у�P   P   Ѓ��у��у��܃�[у�_ڃ�N؃�tك�b���6ރ��⃽�׃�]ރ��׃��ԃ��փ�(Ӄ�Ѓ�9Ѓ��Ƀ�P   P   ̓��ԃ��у��Ѓ�#у�3ڃ��ރ��ڃ��䃽Cك�ۃ�ჽ�܃�I܃��؃��҃�fЃ�TЃ�iӃ�tσ�P   P   �ƃ�Gƃ�ȃ�F̃�ƃ�l̃�!˃��у�ك��׃�u߃�PՃ��݃��΃�Ѓ�ʃ�Ń�Ƀ�dƃ�xŃ�P   P   xŃ��ă��ă��ƃ��ʃ��˃�Pԃ��҃��݃�ރ��⃽\���%܃��ۃ�_փ�C΃�#̓��̃�]ƃ��ƃ�P   P   dƃ�����
ă��ƃ��˃�rӃ��փ�Cヽ�ჽ�䃽�惽V�냽}���Pჽ�⃽�փ��Ճ�Mȃ�]ƃ�P   P   Ƀ��ă��ƃ�9΃�:ǃ��ԃ��փ�k؃��都�ヽ�能}ヽ�僽能�䃽 烽܃�xу��Ճ��̃�P   P   Ń�ʃ�qǃ��ʃ��ǃ�̃��ۃ��ԃ�.烽7샽C�������3냽E��������܃��փ�#̓�P   P   ʃ�7Ƀ��ǃ�LÃ��ǃ��ʃ�у��߃� 能W�샽�􃽘b����샽K��� 烽�⃽C΃�P   P   Ѓ��Ѓ��Ƀ�rɃ�vɃ��σ�Ĩ��փ�䃽�䃽k����
���c����샽�󃽽䃽Pჽ_փ�P   P   �΃�^Ƀ��˃�Bσ��у�
˃�,˃�6у�ڃ��݃�'ꃽQ����$��
���b���E���能}����ۃ�P   P   �݃��у��ȃ��Ã�[ȃ�2ǃ��Ń�ԃ��ك�����+都s能�都���3냽�僽�냽%܃�P   P   PՃ��ԃ�Ƀ��Ƀ�ƃ��Ń�nɃ��̃�Ѓ�Kփ��ヽ�烽s能Q������􃽠���}ヽV\���P   P   u߃�'؃�1Ń�Fʃ��˃��ă�[ǃ�-Ƀ�ă��؃�U݃��ヽ+都'ꃽk򃽇샽C����能�惽�⃽P   P   �׃�]ۃ�UɃ�xǃ�����%������zÃ�/Ń�3̓��؃�Kփ������݃��䃽W7샽�ヽ�䃽ރ�P   P   ك��Ѓ�VÃ�ƃ�������%�廃��Ã�/Ń�ă�Ѓ��ك�ڃ�䃽 能.烽�都�ჽ�݃�P   P   �у�փ�[̃��ʃ�Oă�ǻ������6Ã�廃�zÃ�-Ƀ��̃�ԃ�6у��փ��߃��ԃ�k؃�Cヽ�҃�P   P   !˃�IɃ�mƃ��˃��ƃ�����;�������%����[ǃ�nɃ��Ń�,˃�Ĩ�у��ۃ��փ��փ�Pԃ�P   P   l̃�0у�q˃�>ȃ�UŃ���������ǻ������%����ă��Ń�2ǃ�
˃��σ��ʃ�̃��ԃ�rӃ��˃�P   P   ƃ��ȃ�eσ�]΃��Ƀ�UŃ��ƃ�Oă��������˃�ƃ�[ȃ��у�vɃ��ǃ��ǃ�:ǃ��˃��ʃ�P   P   F̃��ʃ��Ã� ȃ�]΃�>ȃ��˃��ʃ�ƃ�xǃ�Fʃ��Ƀ��Ã�Bσ�rɃ�LÃ��ʃ�9΃��ƃ��ƃ�P   P   ȃ��Ń��ǃ��Ã�eσ�q˃�mƃ�[̃�VÃ�UɃ�1Ń�Ƀ��ȃ��˃��Ƀ��ǃ�qǃ��ƃ�
ă��ă�P   P   Gƃ������Ń��ʃ��ȃ�0у�IɃ�փ��Ѓ�]ۃ�'؃��ԃ��у�^Ƀ��Ѓ�7Ƀ�ʃ��ă������ă�P   P   䧃�����"���b���
ă��Ń�cЃ��փ��σ��փ�ۃ�؃��΃��փ�;σ�1Ń�������$������P   P   ���|���躃�����ƿ���Ń�Hʃ��؃��Ӄ�+݃��҃�%׃��؃�;Ճ��׃�5Ƀ�Sƃ�L������Ӹ��P   P   $���ȴ������ٺ��򻃽�ȃ�t˃�ԃ�ك�}僽�탽�ヽ��僽�ڃ��σ�VЃ���纃����P   P   ����&������ʶ��𺃽����Jփ�Ӄ�⃽�能V����o���냽/݃��փ�lԃ���L���P   P   ��*�������޶��yŃ��ǃ��Ѓ� ׃�k߃��都`냽��������>ꃽ탽܃��փ�VЃ�Sƃ�P   P   1Ń���������I��������ǃ��ǃ��΃��߃��烽������A���
��b����탽/݃��σ�5Ƀ�P   P   ;σ�W���ߵ��h���l�������cσ�k׃��ރ��惽���������������� ��b���>ꃽ�냽�ڃ��׃�P   P   �փ�"ǃ�����s���˺��û��#ȃ�6փ�dԃ�僽b����󃽨�����������
������僽;Ճ�P   P   �΃��Ƀ��ă�6���
�������Ń�$ʃ�˃�7܃� �������|����������A������o���؃�P   P   ؃��ƃ�ȃ���������~�������)ǃ�>ʃ�}׃��Ճ�K⃽�����󃽁���������􃽀ヽ%׃�P   P   ۃ��Ƀ��Ã�����鶃�>�������ÿ������΃�ԃ��Ճ� ���b���������`냽V����탽�҃�P   P   �փ�e΃�wǃ�,Ń�����4�������<����ƃ��ă��΃�}׃�7܃�僽�惽�烽�都�能}僽+݃�P   P   �σ��ă��ƃ��Ń��������������������ƃ����>ʃ�˃�dԃ��ރ��߃�k߃�⃽ك��Ӄ�P   P   �փ��̃��ƃ�l���o���n������T�������<���ÿ��)ǃ�$ʃ�6փ�k׃��΃� ׃�Ӄ�ԃ��؃�P   P   cЃ��ȃ�iŃ�o���ฃ�O���གྷ��������������������Ń�#ȃ�cσ��ǃ��Ѓ�Jփ�t˃�Hʃ�P   P   �Ń�뽃���� ���Ļ�����O���n�������4���>���~������û�������ǃ��ǃ������ȃ��Ń�P   P   
ă�����C������괃�Ļ��ฃ�o�����������鶃�����
���˺��l�������yŃ�𺃽򻃽ƿ��P   P   b������������������ ���o���l����Ń�,Ń���������6���s���h���I���޶��ʶ��ٺ������P   P   "������縃�����C������iŃ��ƃ��ƃ�wǃ��Ã�ȃ��ă�����ߵ�����������������躃�P   P   ������������������뽃��ȃ��̃��ă�e΃��Ƀ��ƃ��Ƀ�"ǃ�W�������*���&���ȴ��|���P   P   ����ԡ�������������|�������L����̃�Aԃ�Ƀ�]փ��ȃ�m���H���ѷ���������{����P   P   �ˣ��Ԝ������S���%������̓�&փ��߃��ヽ!䃽�݃��Ճ�#ʃ��ǃ�6�������ê�����P   P   {���>���n���&�������(����Ƀ�2Ѓ��܃�Zۃ�.���E惽�ۃ�G߃�܃�Ѓ��Ń�K���,���ê��P   P   ���ǫ��
���ݦ�������������e؃��ۃ�A탽e냽M�������V탽~都�߃��փ�����K�������P   P   ��������橃�~������������Ã�<܃�H⃽|탽����Q�����������h能b惽�փ��Ń�6���P   P   ѷ��,���߬��ృ���������Ń��σ�����>能]�������b ��������'���h能�߃�Ѓ��ǃ�P   P   H���l���*���K������R���e��� ʃ��ڃ�ꃽ(����������C��o��������~都܃�#ʃ�P   P   m���͸����������ͣ��"�������a���sՃ��߃��냽��d���u��C����������V탽G߃��Ճ�P   P   �ȃ�u�����������������ұ��ִ��}̓��ك�m߃����� ��d������b ��Q��������ۃ��݃�P   P   ]փ��Ã�_�������+��������������rŃ��Ӄ�rჽ�샽�����􃽣��������M���E惽!䃽P   P   Ƀ������������g������k�������Ǽ��㹃�`˃�rჽm߃��냽(���]������e냽.����ヽP   P   Aԃ���������~���짃��������������������㹃��Ӄ��ك��߃�ꃽ>能|탽A탽Zۃ��߃�P   P   �̃��ƃ�׿������������� ���ݢ��8�������Ǽ��rŃ�}̓�sՃ��ڃ�����H⃽�ۃ��܃�&փ�P   P   L���D������ ������|����������ݢ�������������ִ��a��� ʃ��σ�<܃�e؃�2Ѓ��̓�P   P   ����ظ��e���䥃�����㟃�������� �������k�������ұ������e����Ń��Ã������Ƀ���P   P   |����������������������㟃�|����������������������"���R��������������(���%���P   P   ���׭������k���(�����������������짃�g���+�������ͣ��������������������S���P   P   ��������%���;���k�������䥃� �������~�����������������K���ృ�~���ݦ��&�������P   P   �������R���%�����������e������׿����������_����������*���߬��橃�
���n���Ԝ��P   P   ԡ��é���������׭�����ظ��D����ƃ����������Ã�u���͸��l���,�������ǫ��>���ˣ��P   P   ��������t���n����������$���w����Ã�����Wʃ�Ŀ��}Ã��������������������L���o���P   P   o���򋃽=������.���E�������%ă�Bփ��у�
ჽtރ�փ��ԃ��ă� �������j�������񕃽P   P   L������Ԕ��-������1����Ã�8΃��߃�1能5샽�$냽�烽|ڃ�\σ�V���������������P   P   ���� ���`�������e���Թ�������̓��ރ����������C��������샽kჽ�ʃ���������j���P   P   �������Q���ꝃ�Ġ��ڪ��󿃽�ǃ��僽��������Y��������}�ヽ�ʃ�V�������P   P   �����������p���3���0���$���FЃ��߃�$�\������P����>�����}�kჽ\σ� ���P   P   ����T�������J�������Ū�����|ă�ك�?���"����o���"�����>������샽|ڃ��ă�P   P   ��������𜃽���G�������#�������,ԃ��能�������������"������������烽�ԃ�P   P   }Ã�K���ȣ��������������������ƃ�{ԃ�M都���������o��P��Y��C���$냽փ�P   P   Ŀ��㶃�����㥃�E���0�������穃�����)����݃�������������������������tރ�P   P   Wʃ�tă��������<�������읃�������������σ��݃�M都����"��\����������5샽
ჽP   P   ��������2���3���ݞ������g���>���󞃽�������)���{ԃ��能?���$����1能�у�P   P   �Ã�����*���\���L���|�������=���񜃽󞃽���������ƃ�,ԃ�ك��߃��僽�ރ��߃�Bփ�P   P   w�����������ؠ��0���}���W�������=���>�������穃��������|ă�FЃ��ǃ��̓�8΃�%ă�P   P   $���g���'������A���ӓ������W�������g���읃���������#������$���󿃽�����Ã�����P   P   ��������s���Q���h���	���ӓ��}���|�����������0�����������Ū��0���ڪ��Թ��1���E���P   P   ������ٞ������ɝ��h���A���0���L���ݞ��<���E������G�������3���Ġ��e������.���P   P   n���󘃽�����������Q������ؠ��\���3������㥃�������J���p���ꝃ�����-������P   P   t���I���������ٞ��s���'�������*���2�����������ȣ��𜃽�������Q���`���Ԕ��=���P   P   ��������I���󘃽�������g���������������tă�㶃�K�������T����������� ������򋃽P   P   k���t��Gt��z������G���c�������SÃ�)˃��̓��ȃ���_����������}����y��8y��dp��P   P   dp���m��Zw������򏃽%���b���h���&σ��ރ��܃��܃��ރ�)σ��Ã�X���Q���+��������u��P   P   8y��b|���y������G�������a����΃�sۃ�o񃽜 ��������OFڃ��̃�5���r�����������P   P   �y��(y��Qv��~��2������������҃�:ꃽJ򃽭�����`
��e��:����都҃�]���r���+���P   P   }���⃃�8������ϓ������N���<Ѓ�l0���������!�����
�����惽҃�5���Q���P   P   ����|���J�������L������;���>σ�-能���M���$��5-���2��%��������都�̃�X���P   P   ���픃�����݄��ш������Q����ă�{܃����	���&���3���-��}7��%��
��:���Fڃ��Ã�P   P   _�������s���R�����������會�˴��΃�	/��o��s3���2���-���2�����e��O)σ�P   P   ��Ԥ��铃�����d������Β��Q�������dჽ�������J��s3���3��5-���!��`
�����ރ�P   P   �ȃ�����_���u����|��
�������H���5����Ƀ�5݃��������o���&���$�������������܃�P   P   �̓�ɱ������T���t�����w������ɕ��0���Jʃ�5݃�����/���	��M��������� ���܃�P   P   )˃�u�������䎃�.p���x���v��=s��񉃽X���0����Ƀ�dჽ	�􃽕��0��J�o񃽽ރ�P   P   SÃ�������������}���r��yu��'n�����񉃽ɕ��5�������΃�{܃�-能l:ꃽsۃ�&σ�P   P   ����٥��M�������
q���r��Ze���d��'n��=s������H���Q���˴���ă�>σ�<Ѓ��҃��΃�h���P   P   c���s������������s��Zy���q��Ze��yu���v��w������Β��會�Q���;���N�������a���b���P   P   G���/��������������؀��Zy���r���r���x�����
������������������������������%���P   P   ����%���Q�������쀃�����s��
q���}��.p��t���|��d������ш��L���ϓ��2���G���򏃽P   P   z��3������򄃽��������������������䎃�T���u�������R���݄���������~����������P   P   Gt���z���������Q�����������M��������������_���铃�s�������J���8���Qv���y��Zw��P   P   �t��r|���z��3���%���/���s���٥������u���ɱ������Ԥ������픃�|���⃃�(y��b|���m��P   P   +Y���K��FX���c��x��[����������ʃ�Gȃ��˃�ü��������Z����t���a���R���O��P   P   �O��JK���O��xk��h��畃�l���2��Ӄ��⃽I能N냽����Ӄ�)ă�Q���d����~���j��L��P   P   �R���W��S���i���z�����y���7΃�*탽X���M��u��A�����u能�ȃ�b�������U|���j��P   P   �a��`^���\��cd��.�������j����ԃ���C��� ���0���1��K!������ԃ����������~��P   P   �t��A^���]���_��9v��^������1ك��ꃽV���8��B��FM���D���6�����#ԃ�b���d���P   P   Z���+t��pe���j��cm������"���qɃ���������=��N���W��bT��0O���<�����󃽦ȃ�Q���P   P   ���t���;t���d���u��S������������ꃽW���9��}K��Uc���m���\��0O���6�����u能)ă�P   P   ���.���U��� g���f�����W���e����҃�����P!��yE���Q��7o���m��bT���D��K!������Ӄ�P   P   ü��#���W��Xr���j��]s�������������,������r0��ZM���Q��Uc���W��FM���1��A�����P   P   �˃�`���鈃��j��>j���h��~n��炃�󧃽H˃�_냽o
��r0��yE��}K��N��B���0��u��N냽P   P   Gȃ�䡃�Փ���}���g���b��b��|������5�������_냽���P!���9���=���8��� ��M��I能P   P   �ʃ�ޣ��\����w���e��]Z���V���f��qw������5���H˃�,�������W�����V��C��X����⃽P   P   ���������'v���\���_��?R��K`��>]��qw������󧃽����҃��ꃽ�����ꃽ��*탽�Ӄ�P   P   �'�������}��xg��f���R��PY��K`���f��|��肃�����e�������qɃ�1ك��ԃ�7΃�2�P   P   �������x����n���e���Z���O���R��?R���V��b��~n������W�������"������j���y���l���P   P   [���
��������r��Zk���c���Z��f���_��]Z���b���h��]s�����S�������^����������畃�P   P   x��pu��yu��Wk���j��Zk���e��xg���\���e���g��>j���j���f���u��cm��9v��.����z��h��P   P   �c��md���h���e��Wk���r���n��}��'v���w���}���j��Xr�� g���d���j���_��cd���i��xk��P   P   FX���[��A\���h��yu������x����������\���Փ��鈃�W��U���;t��pe���]���\��S���O��P   P   �K���Y���[��md��pu��
�������'�������ޣ��䡃�`���#���.���t���+t��A^��`^���W��JK��P   P   ���� ���5���J��L[��
y������g��������Ã�&σ��ă�����s������ku��\���J��1���!��P   P   �!���'��x9���:��?U���{��֠����T⃽���� �����ރ�[�������z���O��v<��z9��P   P   1������4��J;���Y��'�������̃�t����&���+���#�������΃�:���܇���U��v<��P   P   �J��?6�� 6��fE��LX�����������ڃ�����)���F��oQ���N���F��W%����ك�Q���܇���O��P   P   \���L��8��)Q���U��}��%����܃�]���6��%U���p��Mu���o��%V��T2��(��ك�:����z��P   P   ku��:\���B��G�� [���w��f����̃����4���X��Q~�����������~��vZ��T2�����΃����P   P   ����d���S��N���O���j������û�����&��U���~��-���r���f����~��%V��W%���[���P   P   s��������O��3O���K��fU���z��
����ჽ����B��br��󐄽s���r��������o���F������ރ�P   P   ���������l��M���I��BK���h������H����샽*(���J��Dz��󐄽-�������Mu���N���#����P   P   �ă�-����j���O���?���;���P���j����������� ��+���J��br���~��Q~���p��oQ���+��� ��P   P   &σ������p��{J���B���/���B�� M���l�����?̃�� ��*(���B��U���X��%U���F���&����P   P   �Ã�U���\���N���D���+���/��cA���M���{����������샽����&��4���6���)�����P   P   ����u���[p��M��+6���%������&��v.���M���l������H����ჽ�􃽀��]�����t�T⃽P   P   g���<���&m���M��JC���&���%���#���&��cA�� M���j������
���û���̃��܃��ڃ��̃���P   P   �������8k��&P��eH���+��O���%������/���B���P���h���z������f���%����������֠��P   P   
y��n���S���Q���?��$2���+���&���%���+���/���;��BK��fU���j���w��}������'����{��P   P   L[��]���O��SO��8N���?��eH��JC��+6���D���B���?���I���K���O�� [���U��LX���Y��?U��P   P   �J���K���K���S��SO���Q��&P���M��M���N��{J���O��M��3O��N��G��)Q��fE��J;���:��P   P   �5���8��=<���K���O���S��8k��&m��[p��\���p���j���l���O���S���B��8�� 6���4��x9��P   P   � ������8���K��]��n�����<���u���U�������-������������d��:\���L��?6������'��P   P   �݂�������y��N:���^����ϟ������mӃ��Ӄ�[΃�}���I���{����]���3��������A삽P   P   A삽�삽����A���@��e��Ǘ���ă��냽;��Z�����:���烽����ߖ���b��F>�����C���P   P   ����?���������`J��Xm������ჽ&
���6��;O��PU��}Q��q2�����0ჽ����n��J�����P   P   �� ��I������&B��sp������惽�&��V��R����������~��wT���!���僽�����n��F>��P   P   �3�������Z���4��a��ӥ��	ヽT-��#o��К������Ą�l���c���kp��J*���僽����b��P   P   �]��1(��������3-���Z�������ჽ�#���o�������Մ��鄽f턽�Є�竄�kp���!��0ჽߖ��P   P   {����O���)��?��%��uR��N}��������tT��;����Ԅ�J�N���T����Є�c���wT���������P   P   I���pd��<��:&��(��h=���a�����a烽Z1���~��𵄽r섽��N���f턽m����~��q2���烽P   P   }���Ku��[H���'��F���(���E��x����������R����������r섽J􄽍鄽�Ą����}Q��:��P   P   [΃������Z���7��������4��Q\�������Ѓ�G
��OR������𵄽�Ԅ��Մ�������PU�����P   P   �Ӄ�|����^���.��H��N
������*���Z��s���Ճ�G
���R���~��;�������К��R���;O��Z��P   P   mӃ�Ζ���[���7��������w���	��V:��h\��s����Ѓ����Z1��tT���o��#o��V���6��;��P   P   ����Ւ��/^��>��w��]��������������V:���Z����������a烽���#��T-���&��&
���냽P   P   ϟ���{���]���0��Y��H�z����邽�����	���*��Q\��x����������ჽ	ヽ惽�ჽ�ă�P   P   ��%d���J��77�����������z�������w�����4���E���a��N}������ӥ���������Ǘ��P   P   �^��V��W@��0�����������H�]������N
������(��h=��uR���Z��a��sp��Xm��e��P   P   N:���-��Q-���)��t��������Y��w�����H�����F��(��%��3-���4��&B��`J���@��P   P   y�����F���$���)��0��77���0��>���7���.���7���'��:&��?�����Z��������A��P   P   ���������F��Q-��W@���J���]��/^���[���^���Z��[H��<���)��������I����������P   P   ������������-��V��%d���{��Ւ��Ζ��|�������Ku��pd���O��1(���� ��?����삽P   P   힂�Š��ʶ��X݂�:��r>���o������4ƃ��߃�P惽܃��ǃ����l���;�����(ڂ�г��R���P   P   R���ך��e���u₽���CP��i���hσ�����)��<���@��{$��j���B΃�ꅃ�M�����ق�R���P   P   г������ܶ���ۂ�,���K��B����냽g3��{f�������������Na���4��L烽Р���E��C���ق�P   P   (ڂ�������[܂����OM��ɲ��
����Q��Ӝ��ʄ� 鄽L焽kƄ�u���2J������M����E����P   P   ����ۂ��Ԃ��ق�I��bK��̢��" ��WP��'���C����!.���������O������Р��M��P   P   �;��� ���낽�肽B��]<��\���}烽M���������8���W���X���7��N������2J��L烽ꅃ�P   P   �l��4&��.�x���x���"��(o��%̃��2�������򄽈4��ie��`}���c���7���u����4��B΃�P   P   ��;M��q��]炽^낽W���N������5����`���Ǆ�)��DU������`}���X�����kƄ�Na��j���P   P   �ǃ�`e��P��b����݂�b����d�������'������Y脽5-��DU��ie���W��!.��L焽����{$��P   P   ܃��{���-����Tڂ�X܂�����P-���x��ރ��<��v���Y脽)���4��8����� 鄽����@��P   P   P惽����<@������ӂ�]Ȃ�Tт�4���>�����������<�������Ǆ������C�ʄ�����<��P   P   �߃������8�������Ȃ�j���Y����Ȃ�.����4������ރ��'���`����������'���Ӝ��{f���)��P   P   4ƃ�D}���@��z���C΂�԰��������͂�.����>���x������5����2��M��WP���Q��g3�����P   P   �����k���1��d���̂��������F�������Ȃ�4��P-���d������%̃�}烽" ��
����냽hσ�P   P   �o���S�����{���҂�����t����������Y���Tт���������N��(o��\���̢��ɲ��B���i���P   P   r>���'��X��h�\₽�ɂ��������԰��j���]Ȃ�X܂�bW��"��]<��bK��OM���K��CP��P   P   :����������킽₽\₽҂��̂�C΂��Ȃ��ӂ�Tڂ��݂�^낽x���B��I�����,�����P   P   X݂��Ⴝ[낽+悽�킽h�{���d��z������������b���]炽x����肽�ق�[܂��ۂ�u₽P   P   ʶ����nۂ�[낽����X������1���@���8��<@���-��P��q��.􂽯낽�Ԃ�����ܶ��e���P   P   Š��Բ�����Ⴝ����'���S���k��D}�����������{��`e��;M��4&��� ���ۂ�������ך��P   P   r;��N;���a��t����Ƃ�����\��J���A̓�Q냽����탽�ă�"����U�����Ă�����^��<��P   P   <��p>��(e�������т��,��y���W؃����]���r��u��Z�����'փ�L���&���̂�揂��`��P   P   �^��A���`������yق�D��w�������f��ɴ���焽����6ℽ0���Ka������v����<���ӂ�揂�P   P   ����i��k��T���'т��>��졃���������򄽦9���`��6[��;���񄽮���K��۞���<���̂�P   P   Ă�W���t��Ҏ��Ƃ�"(��4���B��W�������v��q����Ņ�崅�3s��Z��.���K��v���&��P   P   ���)Ȃ�T�������%Â�G��;�����������������+ㅽ7��	���慽ш��Z����������L���P   P   �U���낽𳂽��������ꂽW���Ӄ�-b����p���ⅽv!���5������慽3s����Ka��'փ�P   P   "������˂���������(ɂ�����������񴄽K6��]���&
��!0���5��	��崅�;��0������P   P   �ă��[���������������������3V���Ń�yT������W��MŅ�&
��v!��7���Ņ�6[��6ℽZ��P   P   탽�k��=��d�������U���-�������*k���ヽs���W��]����ⅽ+ㅽq����`������u��P   P   ����c������{���0���Vt���������u������y탽s������K6���p������v���9���焽�r��P   P   Q냽$���K'��������c���a��W���K���"�������ヽyT��񴄽���������ɴ��]��P   P   A̓��o��a��N��������[��MG���X���|��K���u��*k���Ń����-b������W��������f�����P   P   J����Y���
���z���a���G���H���X��W����������3V�������Ӄ�����B��������W؃�P   P   �\��(�������������ne���E���G��MG���a������-����������W��;���4���졃�w���y���P   P   ���񂽊҂�J���瓂��v��ne��a���[���c��Vt��U������(ɂ��ꂽG��"(���>��D���,��P   P   �Ƃ��ʂ������������瓂�����z����������0������������������%Â�Ƃ�'т�yق��т�P   P   t������k���0�������J��������N�����{���d�������������������Ҏ��T�����������P   P   �a���o��.t��k��������҂�����
��a��K'�����=�������˂�𳂽T���t��k���`��(e��P   P   N;��H���o������ʂ��(���Y���o��$���c����k���[�����낽)Ȃ�W����i��A��p>��P   P   ����º��^���R/��}���Ⴝ$I������n能���������ჽ	���fG���ق��z��`&���ၽ+���P   P   +���]����؁��������r����w��^�G\�������Ǆ����螄��Y��s탽�r�����������ց�P   P   �ၽX΁��ށ����@���
�������7��3������^��]y��-Y�����Y����3������	��΋�����P   P   `&���������a'�������������_T��儽�q���څ�x�����Gۅ��k���焽/L�������	������P   P   �z���0������3���w���������	N���󄽘���'���y��򘆽Oz��%���������/L�������P   P   �ق�l���.���.���l���؂�.v��k6��1ㄽ�����>��|�����솽W����B�������焽�3���r��P   P   fG������_��?��\[��/�A���샽����l��C"��|���t���1�����W���%���k��Y���s탽P   P   	�������8��A��>���~��������T������څ��w��,�,���1���솽Oz��Gۅ�����Y��P   P   �ჽ$.������M��E.��Q��§���*��N⃽V����Y�����8���,t���򘆽���-Y��螄�P   P   ����b��0˂�%`��e%���!���^��ł�[^�����u����s������w��|���|����y��x��]y�����P   P   ��
p���؂�	`��O������K��;\��gԂ��h��E��u����Y���څ�C"���>��'���څ��^���Ǆ�P   P   ���sp���₽�r�����t䁽<䁽
���m���ق��h�����V�������l�����������q��������P   P   n能2f���݂��p�����Oρ������΁����m��gԂ�[^��N⃽�T�����1ㄽ��儽3���G\��P   P   �����2���΂��e�����Ӂ�ǵ�������΁�
��;\��ł��*������샽k6��	N��_T���7��^�P   P   $I���������c������災�Ł�ǵ������<䁽K���^��§����A��.v���������������w��P   P   �Ⴝ�Ƃ� ���X���(�����災Ӂ�Oρ�t䁽�����!��Q���~��/��؂�������
��r���P   P   }���t��@a���I���5���(��������������O��e%��E.��>��\[���l���w������@�������P   P   R/���7���:���D���I��X��c���e���p���r��	`��%`���M��A��?���.���3��a'��������P   P   ^���K�������:��@a�� �������΂��݂��₽�؂�/˂����8���_���.���������ށ��؁�P   P   º���Ӂ�K����7���t���Ƃ������2��2f��sp��
p���b��$.���������l���0������X΁�]���P   P   �瀽V��(B��n����������
������Z����7��jT��	3������D�����b���������n@�����P   P   �����m;�������#���Ȃ�d��
����������<��~:��M���㚄����\����5��Ҝ��7��P   P   n@��n(���?����������Ђ����j_�����񮅽���1��I��{�������\��^���|Ȃ�>��Ҝ��P   P   ���H��8K������n��Cт�񹃽=���u���6��򺆽����b���;����4���p��/���w���|Ȃ�5��P   P   �������C{��v����������������鈅��x���)��:���|Ƈ�����*���w���}��/���^�����P   P   b����끽%���Ψ����Z���;X��^���p��}y��N��󇽠F��~I��y����Q���w���p���\���\��P   P   ���R��݁�C���ځ��S��Z��;��J��W1���(��&򇽷u������|��y����*���4�������P   P   D���＂�"��ʁ�h΁�W��D���v������K���2���=����G��ɝ�����~I�����;���{���㚄�P   P   ������K��ځ�y���a؁�wE������Y탽�������������G���u���F��|Ƈ�b���I��M���P   P   	3��H���{��J큽ݢ��ខ��恽�{��=��W.��)3��|%������=���&��:��������1��~:��P   P   jT���i��Ꞃ�����܋��Gl��������������\��uO��)3����2����(��N���)��򺆽���<��P   P   �7��4l��������U����G���H��e{��w���K����\��W.������K���W1��}y���x���6��񮅽���P   P   Z����H��|������i��� =�����59��F���w�������=��Y탽���J���p��鈅�u���������P   P   �������e���|�����	=��p
�����59��e{�������{������v���<��^������=���j_��
��P   P   
�����cU��?�H���_L��9#��p
������H������恽wE��D���Z��;X������񹃽���d��P   P   �����^���&��J偽����6u��_L��	=�� =���G��Gl��ខ�a؁�W���S��Z�����Cт��Ђ��Ȃ�P   P   �������遽=ց���������H������i���U���܋��ݢ��y���h΁�ځ��򁽺��n������#��P   P   n���i�������5Ɓ�=ց�J偽?�|������������J큽ځ�ʁ�C���Ψ��v���������������P   P   (B���Q��X�������遽�&��cU��e���|������Ꞃ��{��K��"��݁�%���C{��8K���?��m;��P   P   V��v)���Q��i��������^���������H��4l���i��H����＂��R���끽����H��n(����P   P   *������f���‽����fC��z���?����"���z��D���'v����������ꂽ�<��Ut��_ۀ�/^�����P   P   ����
���O���ۀ�����r���l���L��� ��𞅽<ׅ�4ۅ�ƕ�������D��f��i��i���mـ�3J��P   P   /^���2���`��$ۀ�ꝁ�ԗ��Z���*�����������g���+�����j�������'���������阁�mـ�P   P   _ۀ�>���X����ހ����S���U���m愽.���(��+�Z���V��f)��:%���ㄽ������i���P   P   Ut��<瀽�����〽$y���k��S����脽%S���������z2���l���2��������S���ㄽ���i��P   P   �<��k��}�C��i��&=��=b��۰���&���|��?�������������q����������:%��'���f��P   P   �ꂽPぽ9@��|���R@���ف��낽�@������D%������٠��]P������~N��q������f)�������D��P   P   �����d��ی�������������a��E������{��:臽�-�����)�����������2��j�������P   P   ���EႽ؁��,��T����)��&ց�{ق����s���N���O��/j�����]P������l���V�����ƕ��P   P   'v���(��\��J@���Ӏ�aЀ�:������!��Ki��Ѕ��%���O���-��٠������z2���Z���+��4ۅ�P   P   D����Y���7��2W��{ɀ������ɀ�6L���)��0S�����Ѕ�N��:臽����?������+g��<ׅ�P   P   �z��]]���L���\��ؾ���a���\��n���MR��C��0S��Ki��s����{��D%���|�������(������𞅽P   P   �"���.���9��9`�������K�����|E��<���MR���)���!������򄽞����&��%S��.������� ��P   P   ?����炽���-[���À�-L��1��Z��|E��n���6L�����{ق�E����@��۰���脽m愽*����L��P   P   z����p���䁽�M���р��i��=#��1������\���ɀ�:��&ց��a���낽=b��S���U���Z����l��P   P   fC����������7���ހ�홀��i��-L���K���a������aЀ��)�������ف�&=���k��S���ԗ��r��P   P   �����u���P���$��3 ���ހ��р��À�����ؾ��{ɀ��Ӏ�T������R@���i��$y�����ꝁ�����P   P   �‽q�����a���$���7���M��-[��8`���\��2W��J@���,�����|���C��〽�ހ�$ۀ��ۀ�P   P   �f��؎��<��������P�������䁽����9���L���7��\��؁�ی��9@��}󀽃���X����`���O��P   P   ���u6��؎��q񀽱u������p���炽�.��]]���Y���(��EႽ�d��Pぽk��<瀽>����2���
��P   P   rK}�ɗ}�D}~�����À�����|���ӛ��(^���܄�c��ۄ��T������)���N����������c~���}�P   P   ��}��}�-]~�w���‽���jE�����ڏ���W��vÆ�6Æ�aR�������w���8�������ۀ�#���Q~�P   P   c~���}�g~�ۭ�;〽N/��ҭ��/��̍�������W������=T��a������'��ȣ��g,��!Ӏ�#��P   P   ���:�~���~�����ހ��*��c̃� ����(������n���wF���>��+�������&��z���6Ã�g,���ۀ�P   P   ����V���0�C������I�����������_h��U$�������m��T����o������?���l��z���ȣ������P   P   N�������>���������렁�n:���!�� '��H��#ފ��������ػ������ߊ�?���&���'���8��P   P   )����E��`�����a���B��_���Wr�������׌����� ��y��h
���������������w��P   P   ���� � Ā�1���&�����큽����T���e�������Vj�������t��y��ػ���o��+���a�������P   P   �T��A����.���P��E���M���&��Ղ���O��wC��J��V2���������� ������T����>��=T��aR��P   P   ۄ����@���Pr��y��3���m���w�������Ʉ��������V2��Vj���������m��wF������6Æ�P   P   c��e@��ں������ϐ����|�恀�����(1��2����J������׌��#ފ�����n����W��vÆ�P   P   �܄��@��ԁ�Ӟ��i�)�~�Q�~��^���������(1���Ʉ�wC��e������H��U$�����������W��P   P   (^�����,���'���;q�W;~�5�}��/~�FR��������������O��T����� '��_h���(��̍��ڏ��P   P   ԛ��q���،��~����x��D~�ׯ}��}��/~��^�恀��w��Ղ������Wr���!������ ���/�����P   P   |��� ���8�����y����~�\�}�ׯ}�5�}�Q�~��|��m���&���큽_���n:������c̃�ҭ��jE��P   P   ����HS��#ր��b����L#���~��D~�W;~�)�~���3���M�����B��렁�I����*��N/�����P   P   �À������n���>��%����y���x�;q�i�ϐ�y��E���&��a�����������ހ�;〽�‽P   P   ���������"���>���b�����~���'���Ӟ������Pr���P��1��������C�����ۭ�w��P   P   D}~�w�~�\K����n��#ր��8��،��,���ԁ�ں��@����.�� Ā�`��>���0���~�g~�-]~�P   P   ɗ}���}�w�~��������HS����q�������@��e@�����A��� ��E������V��:�~���}��}�P   P   �yy�3z�`={�0}��|����x��Ӻ��	���JX��ĕ��CS��ᬄ�����j��-���_���|��*{�J	z�P   P   J	z��z�{���|�J��Q����8���儽yn��9t��H��x��bo���c��\ڄ�)���u��T����|�n{�P   P   �*{�y�z��.{���|�������rÃ��̅�b���,Q���K�������H��K��Z����ǅ���������q����|�P   P   ��|�ԗ{�8�{�c�|�������j߃�yD�����������#��z)����!��r���o����?���׃�����T��P   P   �_��}��l|�}�!f�x��t���k;�������S���J��E������b���}J���U��E؈��?�������u��P   P   -����~��K}�F}���~�j����'��ܿ������^V��R����y��#y��"z��My������U��o����ǅ�)��P   P   j���k���E~�f�}�G@~��j��m_��3ׄ���������A���x��tꐽ Y���My��}J��r���Z���\ڄ�P   P   �����f��?�%�}�^�}�uv��_��\����X���<�����[���Ru�� Q�� Y��"z��b����!��K���c��P   P   ᬄ�/���K��Y#~�':}��~�g=���#������[��]<���������Ru��tꐽ#y�����)����H��bo��P   P   CS��ق��Ā���~���|���|�"n~�����.Ă��=���󇽆�������[����x���y��E���z����x��P   P   ĕ���0��1��?�~���|���{�!�|�H�~�H��"��������]<������A��R����J���#���K��H��P   P   JX���0��L(���~���|�WA{�D{�|r|�5�~����"���=���[���<�����^V���S������,Q��:t��P   P   	����������N�~���|���z�bz�I�z��^|�5�~�H��.Ă�����X������������������b���yn��P   P   Ӻ��T?���р�1�~�X�|��{��z���y�I�z�|r|�H�~������#��\���3ׄ�ܿ��k;��yD���̅��儽P   P   x���t��\Z���~���|��X{��wz��z�bz�D{�!�|�"n~�g=���_��m_���'��t���j߃�rÃ��8��P   P   ���M�����T~��}�W|��X{��{���z�WA{���{���|��~�uv��j��j���x��������Q���P   P   �|�6�~��u~�5�}�|l}��}���|�X�|���|���|���|���|�':}�^�}�G@~���~�!f�������J��P   P   0}�9}�rv}�.�}�5�}��T~��~�1�~�N�~��~�?�~��~�Y#~�%�}�f�}�F}�}�d�|���|���|�P   P   `={��{�U�|�rv}��u~���\Z���р����L(��1���Ā��K��?��E~��K}��l|�9�{��.{�{�P   P   3z���z��{�9}�6�~�L���t��T?�������0���0��ق�/���f���k����~��}�՗{�y�z��z�P   P   �u��mu�w�v��wy�ƒ|�� ������	����+������f��a��� ��觃��恽N���k|��Ny�|�v�$Yu�P   P   $Yu��Zu�*�v�Yfy���|�o���%��w���z��G��׉��ԉ��	��'q��Xg��������e�|�|Oy�=�v�P   P   |�v�Tv�2�v�Ney�]7}�d���Ӄ�K���di��󕋽	���w��+������`��*���Ƀ�����.}�|Oy�P   P   �Ny�|w�yw��Xy���|�k
��t��kd��S���4y�����S�������{���wx��S����\�������e�|�P   P   �k|��ry�XOx��ny�.p|�̞��O̓��Z�����Ç���Q��1���˓��.���O����������\��Ƀ�����P   P   N����{���y�ۓy�.�{�������6���]��������瑽q��o���<Õ��t���ꑽ����S���*�����P   P   �恽�r~��{�,�y��{�pa~��݁�H[��U���i��
H���n���z���4������t���O��wx���`��Xg��P   P   觃������|�az�gz���|��z������zY��7z�����������4���4��<Õ��.��{������'q��P   P   � ������/;~�H�z�V�y���z�O~���������򈽖�n���X�������z��o����˓�����+���	��P   P   a��c���8v�5c{��Vy�0Oy��F{�HS������������W��n������n��q��1��S����w���ԉ�P   P   �f��j���%����{���x�jx�2�x���{���~���EG����������
H���瑽�Q�����	��׉�P   P   ���"��(W��y|���x�.w�'w��x���{��<��~���������7z���i������Ç��4y��󕋽G��P   P   �+�������.���|���x�&�v�B�u���v���x���{���������zY��U��]������S���di���z��P   P   	����с�W����{�E�x���v�Ԙu���u���v��x���{�HS���������H[��6����Z��ld��K���w��P   P   ����C����q~���{��&y��1w�%�u�Ԙu�B�u�'w�2�x��F{�O~��z���݁����O̓�t���Ӄ�%��P   P   � ��v�~���|�V{���y��6x��1w���v�&�v�.w�jx�0Oy���z���|�pa~����̞��k
��d��o���P   P   ƒ|�|��\{� �z���y���y��&y�D�x���x���x���x��Vy�V�y�gz��{�.�{�/p|���|�^7}���|�P   P   �wy���y�R�y��#z� �z�V{���{���{��|�x|���{�5c{�H�z�az�,�y�ۓy��ny��Xy�Ney�Zfy�P   P   w�v�{�w�t}x�R�y��\{���|��q~�W���.��(W���%��8v�/;~��|��{���y�XOx�yw�2�v�*�v�P   P   �mu�.$v�{�w���y�|�v�~�C����с�����"��j��b������������r~���{��ry�|w�Tv��Zu�P   P   \n�]	o��<q���t���x�8�}������냽����F'��	���� ���ʅ��؃�jd���}���x�qt��q�]o�P   P   ]o�M�n���p�^_t��ey�\��T��O��b!��aC���e���h��9�����i<��
���q\��By�vEt���p�P   P   �q���o�_q��Vt��py�I#������9���>͋�����V鐽㖑�Vᐽ|׎��ċ�9򇽉샽���ay�vEt�P   P   qt���q���q�Vnt��Ry�Y���S�����~�����Ǝ��s/���-��Z������&z��툽>Q������By�P   P   ��x�1ut�B
s�4wt�*�x�}W��都�9��L����������ɞ����
쒽j��툽�샽q\�P   P   �}���w�5�t���t���w�0�}�b悽P釽�o��kⒽ�ї��k��c���_���u��Yח�
쒽&z��9�
���P   P   jd���i{�8�v��"u��v�MM{�^���(�������{����c���]��oy���`���u��������ċ�i<��P   P   �؃��
�c�x�#�u�w�u�H�x���~�b�����������q������,T��	t��py���_��ɞ��Z���|׎����P   P   �ʅ��$����z�Liv���t�]Kv���z����%������!���,��ɀ��,T���]��c������-��Vᐽ9��P   P   � ���Q��6�|�ow��/t��t�q�v� �|�W-������|?��Qs��,�������c���k������s/��㖑��h��P   P   	���������}���w�T�s�-]r�ȭs��w�K�}��΂��d��|?��!����q����ї���Ǝ��V鐽�e��P   P   F'��g����`~�� x�E�s�Lq�&0q��ms���w�~��΂�������������{��kⒽL��������aC��P   P   ����W^���}��.x�ʃs�P�p��o���p��Vs���w�L�}�W-��%�����������o��9���~��?͋�c!��P   P   �냽25����|���w�^�s���p��(o�(o���p��ms��w� �|����c����(��P釽���9���O��P   P   ���?�3{�Vw�T�s��nq���o��(o��o�&0q�ȭs�q�v���z���~�^��b悽�都�S������U��P   P   8�}���{�y�'�v�?tt�̑r��nq���p�P�p�Lq�-]r��t�]Kv�H�x�MM{�0�}�~W�Y��I#��\��P   P   ��x�5�w��w���u��5u�?tt�S�s�^�s�ʃs�E�s�T�s��/t���t�w�u��v���w�*�x��Ry��py��ey�P   P   ��t��t�u�Nsu���u�&�v�Vw���w��.x�� x���w�nw�Liv�#�u��"u���t�4wt�Vnt��Vt�^_t�P   P   �<q���q��Fs�u��w�y�3{���|��}��`~���}�6�|���z�c�x�8�v�5�t�B
s���q�_q���p�P   P   ]	o�� p���q��t�5�w���{��?�25��W^��g��������Q���$���
��i{���w�1ut���q���o�M�n�P   P   :�e�Q�f�f|i�V�m���s�C]z�7�������І������<��ʖ�����#�p���x z��ys� �m��Ti���f�P   P   ��f���f��(i���m���t��|��ׂ�/S��O]��&T��T��쏽-J��'N���;��Â�L�|��\t���m��i�P   P   �Ti���g�Dai��m���t���}��G���Չ�Z��W{���W��xf��lP��s��.	��fȉ�
5����}�Z�t���m�P   P    �m��Uj��]j��m�nt���}�沄��-��]���jW����������.���1���Q�������'��������}��\t�P   P   �ys���m�l�\�m��ns���|�n/���#��dp��d��������S�����$���h���v���'��
5��L�|�P   P   x z��-r��,n��#n�G r��
z����������{��RX��"Q��:���B���Ř��g����_���h������fȉ�Â�P   P   p����*w���p���n�D�p��w�2~���"��i鎽o5��/	��(�������|����g����$��Q��/	���;��P   P   #󃽈|�?�s�>�o�xto�"�s�r�{�v̓��&��9J���w���Ԣ�W���}n���|��Ř����1���	s��'N��P   P   ���x0��ɖv��~p�kkn�N_p��hv��	���������B���Ɲ�1��X������B����S��.���lP��.J��P   P   ʖ��D큽Cy��q�܋m�qm��Yq�}�x�[����Y��Q����1���Ɲ��Ԣ�(���:���������xf���쏽P   P   �<��N܂���z��Rr��m�"Pk�J�l��	r�;Wz�1�������Q���B���w��/	��"Q����������W��U�P   P   �����܂��F{�D�r�w�l�h�i� �i�یl��pr���z�1����Y�����9J��o5��RX��d��jW��X{��&T��P   P   �І�����z���r���l���h�h�g���h���l��pr�;Wz�[��������&��i鎽�{��dp��^���Z��O]��P   P   ����H���?y�izr��l�$i���f���f���h�یl��	r�}�x��	��v̓��"�������#���-���Չ�/S��P   P   7����V|�q�v���q�	Tm���i�2�g���f�g�g� �i�J�l��Yq��hv�s�{�2~������n/��沄��G���ׂ�P   P   C]z��qw�Dt���p���m��k���i�$i���h�h�i�"Pk�qm�N_p�"�s��w��
z���|���}���}��|�P   P   ��s��|r�Zq���o���n���m�	Tm��l���l�w�l��m�܋m�kkn�xto�E�p�H r��ns�nt���t���t�P   P   V�m�n��{n�9o���o���p���q�izr���r�D�r��Rr��q��~p�>�o���n��#n�\�m��m��m���m�P   P   f|i��j�Ul��{n�Zq�Dt�p�v��?y���z��F{���z�By�ɖv�?�s���p��,n�l��]j�Dai��(i�P   P   Q�f��h��j�n��|r��qw��V|��H�����܂�N܂�C큽x0���|��*w��-r���m��Uj���g���f�P   P   FqZ�K�[�J6_�i0e�G�l�~�u����(X��6#����������0���F���4���=�^�u�W�l�l�d�o_���[�P   P   ��[�o�[�߳^��e�T�m���x������䈽�x������� ��+��������e��8ˈ�����y�x�l�m���d��^�P   P   o_�{)]�2_���d��Vn���z�����@\��y��������������L噽N����P��������z�>n���d�P   P   l�d��b`��X`�c�d��m�[�z�?�����[;��Bi��Zƥ��%���%������?f��J7�� ��F:����z�l�m�P   P   W�l��e�#bb�Ne�əl�q�x��~��f��rg���d��ժ�녰��o��S����ت�	s���l�� ������y�x�P   P   _�u���j��]e�jMe���j���u����F3��j��gZ��m����q��᳸�<���@�����	s��K7���P������P   P   �=��wq�g�h��f���h�fLq�W�~�����T���7��ٯ���a��𺽖I��Z��@���ت�?f��N���8ˈ�P   P   �4��5'x�\�l�*"g�g�O�l�j�w����`*�����r���iU��ɞ���A���I��<���S�������L噽�e��P   P   F���1~���p�Vmh���e��@h�/{p�O�}��ɇ��]���ɝ�1䨽�<��ɞ���᳸��o���%���������P   P   0���nf��Kt�%�i�P~d�yd�v�i���s����ZJ��e����.��1䨽jU���a���q��녰��%�����+���P   P   ���������Ov�F�j��c�͂a���c�]�j���u��O��f.��e����ɝ�s���ٯ��n���ժ�Zƥ����� ��P   P   �������2*w��k�$�c�st_��c_�Mgc��Ck�7�v��O��ZJ���]������7��hZ���d��Ci���򙽮���P   P   6#��wz���tv���k�©c�ߊ^���\��Y^��<c��Ck���u�����ɇ�`*��T��j��rg��\;��z����x��P   P   (X���}~��Bt�{(k���c�Q�^�1\�t�[��Y^�Mgc�]�j���s�P�}��������F3��f�����@\���䈽P   P   ����xx��q�sj�Ad��_���\�1\���\��c_���c�v�i�/{p�j�w�X�~�����~��?����������P   P   ~�u�i�q��Bm���h���d���a��_�Q�^�ߊ^�st_�͂a�yd��@h�O�l�gLq���u�q�x�[�z���z���x�P   P   H�l��Uk��ai���g��f���d�Ad���c�©c�$�c��c�P~d���e�g���h���j�əl��m��Vn�U�m�P   P   i0e��de���e�I�f���g���h�sj�z(k���k��k�F�j�$�i�Vmh�*"g��f�jMe�Ne�c�d���d��e�P   P   K6_���`�a�b���e��ai��Bm��q��Bt��tv�2*w��Ov�Jt���p�\�l�g�h��]e�#bb��X`�2_�߳^�P   P   K�[��O]���`��de��Uk�i�q��xx��}~�vz���������nf���1~�5'x��wq���j��e��b`�{)]�o�[�P   P   ةK�.=M�O�Q���Y���c���o�{�|�&���ȉ�7U�������D������k��1R|��Zo�XSc�FHY��Q�(M�P   P   (M��"M��YQ�:mY�0e��t��Q��Hފ����	����𛽯훽!�������Ê�:/��u�s�$e��FY��?Q�P   P   �Q��:O���Q�;ZY���e��Av��������1��o����O$��;��Z���%��噏��鄽/v� ve��FY�P   P   FHY��_S�\S�qJY��d�i"v�S�R���>������?���S��CS��i>������6��UT���/v�$e�P   P   XSc��NY��V�>HY��<c���s��ք��=���꠽c`��^ܻ�zaĽ�nǽ�hĽ�黽�r�����UT���鄽u�s�P   P   �Zo���`��Y�v�Y�C�`�)'o�2	��\o����H�������hʽ�ѽ�
ѽۀʽ?����r���6��噏�:/��P   P   2R|��i�Dp^�̔Z��K^��bi���{�r����♽�˪�����Nʽ�VԽؽkiԽۀʽ�黽����%��Ê�P   P   �k����r��c�k�[���[��_c��;r��!��9:��'����䳽�Ľ@�нE�׽ؽ�
ѽ�hĽi>��[������P   P   �����z�$�h�!�]��Z�'�]��jh�YUz�nN��c0�����}$ǽ@�н�VԽ�ѽ�nǽCS��;��"���P   P   �D��最�]m���_�;�X�m�X�c_���l��7���Ҍ�q��o���}�Ľ�Nʽ�hʽzaĽ�S��O$���훽P   P   �����[���rp��[a�I#X�=�T��W���`��o��ꁽa��q������䳽�������_ܻ��?������P   P   7U���h���q��Bb���W��qR��TR��}W�e�a���p��ꁽ�Ҍ�d0��'����˪�H��c`�����p��
���P   P   ȉ�����-�p��[b���W��7Q��O���P��1W�e�a��o��7��nN��::���♽���꠽�>��1�����P   P   &���@{��m���a��X��JQ���M���M���P��}W���`���l�YUz��!��r���\o���=���R�����Hފ�P   P   |�|�	s��@i�"!`��sX���R��>O���M��O��TR��W�c_��jh��;r���{�3	���ք�S�����Q��P   P   ��o�<j�md��_^��aY��KU���R��JQ��7Q��qR�=�T�m�X�(�]��_c��bi�*'o�«s�j"v��Av��t�P   P   ��c��Va���^�h�\�һZ��aY��sX��X���W���W�I#X�:�X��Z���[��K^�C�`��<c��d���e�0e�P   P   ��Y���Y��CZ�01[�h�\��_^�"!`���a��[b��Bb��[a���_�!�]�k�[�̔Z�v�Y�>HY�qJY�<ZY�;mY�P   P   O�Q�;�S��tV��CZ���^�md��@i��m�-�p��q��rp�]m�$�h��c�Dp^��Y��V�\S���Q��YQ�P   P   .=M��dO�;�S���Y��Va�<j�	s�@{������h���[��圀���z���r��i���`��NY��_S��:O��"M�P   P   Є8�"�:���@�'7J��oW��Ag��x��Є����c�������됽\���)���L?x�_�f��W�G�I��J@���:�P   P   ��:�V�:��?�m9J�,�Y��m�����N���!h���頽m���2����֠��H��wb��������l��ZY�J��?�P   P   �J@��=��]@��J��DZ��p�"g���:��� ��֯������˻�d����˯�`����%��1\��`�o�0Z�J�P   P   G�I�RIB��EB���I�iWY�0�o������◽�/��R���tRɽ�ѽ�ѽUɽ�����1���痽=���`�o��ZY�P   P   �W�B
J���E���I�a�V���l��6��:˗�+����½�Խ0�Ὧ����z�ԽZ½�֬��痽1\����l�P   P   _�f���S��mJ��eJ�z�S��f�g���哽墳������ؽs^�J������-��ٽZ½�1���%������P   P   L?x��x_���P��PK��MP�_�n�w���|����3�� �Խ�8�1,��ux ��V��-��{�Խ����`���wb��P   P   )���yVk��bW��NM��.M�)W��j��<��|Η��A����Ƚ�}�����g �ux ������Uɽ�˯��H��P   P   \���w[v��-^���O���J�(ZO�$�]�~u�n���6�����_cн�2����1,��K�����潑ѽe����֠�P   P   �됽P�~�(<d��AR�+3I�rI���Q��qc��}��C��SϤ����_cн�}Ὕ8�t^�1���ѽ�˻�3���P   P   ���j؁��Vh�	zT�fH��ID�H���S��Tg��>��TϤ� �����Ƚ�Խ��ؽ�ԽuRɽ����n���P   P   d����災�i��U��H�A�W�@���G�[�T�S�h��>���C���6���A���3�������½S���֯��頽P   P   ���9���h�S�U��<H�`�?��<�Hi?���G�[�T��Tg��}�n��|Η�}���墳+����/��� ��!h��P   P   �Є�_�v���d� �T��OH���?�r{;�!T;�Hi?���G���S��qc�u��<�����哽;˗��◽�:��N���P   P   �x���k��^���R���H�r�A��#=�r{;��<�W�@�H���Q�$�]��j�o�w�g���6������#g������P   P   �Ag�5�_�)�W��;P�d�I�z�D�r�A���?�`�?�A��ID�rI�(ZO�)W�_��f���l�1�o��p��m�P   P   �oW��rT��Q��M�sK�c�I���H��OH��<H��H�fH�*3I���J��.M��MP�{�S�b�V�jWY��DZ�-�Y�P   P   '7J��~J�B�J��L��M��;P���R���T�S�U��U�zT��AR���O��NM��PK��eJ���I���I��J�m9J�P   P   ��@�u�B�}-F�B�J��Q�(�W��^���d���h��i��Vh�'<d��-^��bW���P��mJ���E��EB��]@��?�P   P   "�:��R=�t�B��~J��rT�4�_���k�^�v�9��災j؁�O�~�w[v�xVk��x_���S�B
J�RIB��=�V�:�P   P   �{ ���"��O*�^�6��*G�d�[��r����8����}���藽Fj��Ƅ������$r�=[���F�76��*���"�P   P   ��"�d�"��^)�8u6���I�;c�򦀽�����㟽����5���)����㫽�ş��������b�p�I�!J6��P)�P   P   �*��&��*�|P6�Q�J�ׄg����� �����B���&�ν��ӽ�ν������;������{g���J� J6�P   P   76��r,��k,�@!6���I�xKg��\���6��@���XMӽP�-��2���V轢Pӽ�����H��Bl��{g�p�I�P   P   ��F��6��N0���5���F���b�*p�����:6���ݽa@�����~_����'k��Pݽ�p���H�������b�P   P   =[��B��_6��C6��SB�U�Z��1�������*����ܽI ��6�L��U���T�Kx �Pݽ����<�����P   P   $r��FQ���=�!�7���=�N�P��Dq�K���e��W�ҽ������S��;!�my��T�(k���Pӽ������P   P   ������`��F�f:���9��AF�G$`�5����������j�罏=�|��B$!��;!�U������V�����ş�P   P   Ƅ��W�o�}�O��*=���6���<��+O�k�n�?�������ͽpA��
�|���S�L��_�2�� �ν�㫽P   P   Gj��s.{���W�n�@�t5��4�� @�@�V���y�%������(yҽpA�=����6����-����ӽ*���P   P   �藽Ҁ�a[]�S�C�SS4��6/�	�3�+�B�p\�m���������ͽj�����I �b@��P�'�ν6���P   P   �}��ڀ�Us_�fE�D4�Vd+�)'+��[3�H^D���]�m��&�����������X�ҽ��ܽ�ݽZMӽC�������P   P   9����s{�I�]��E��*4���)���%�)0)�wS3�H^D�p\���y�@�����e���*��;6��A�������㟽P   P   ���dp��EX�v�C�^P4���)�y$��Q$�)0)��[3�+�B�@�V�k�n�5���L����������6��� ������P   P   �r��~a��P�+7A�$�4���+�2V&�y$���%�)'+�	�3�� @��+O�G$`��Dq��1��*p���\�����󦀽P   P   e�[�C�Q�9oG���=���5��/���+���)���)�Vd+��6/��4���<��AF�O�P�V�Z���b�zKg�لg�	;c�P   P   �*G�*C�p�>���:�z�7���5�#�4�]P4��*4�D4�SS4�t5���6���9���=��SB���F���I�R�J���I�P   P   _�6���6��7���8���:���=�*7A�u�C��E�fE�R�C�n�@��*=�f:�!�7��C6���5�A!6�}P6�8u6�P   P   �O*��,���0��7�o�>�9oG��P��EX�H�]�Ts_�`[]���W�}�O��F���=��_6��N0��k,��*��^)�P   P   ��"�I&��,���6�*C�C�Q��~a�cp��s{�ڀ�Ҁ�r.{�V�o���`��FQ��B��6��r,��&�d�"�P   P   `"��������ޜ1��K�l�i����(���b���r�������v��܃�!i��dK� =1��w�J�����P   P   ���l����
�^5��U��3}�z[��Ϊ�������ĽS�Ľ�غ����� 2��p�|�ˡU�3.5�B����P   P   J��n����Q��ـ6��S[��[���n��Cs����ڽ��f���а�m�ڽi]���d���T���U[���6�B��P   P   �w��p�Og��]�+�4�X[�ָ��v����ν@���m#���D��z'�M���B�νݨ��݇��U[�3.5�P   P    =1���P�����0�� U����Xy���2Խ_V�����*��X1���*�y�����Y�Խݨ��T��ˡU�P   P   �dK���+�0���T��F+�w�J���{�Ԡ�yBν.�8����7�N�F�"�F��8�<#����C�ν�d��q�|�P   P   !i�v�>�G�%���l�%�i�=���g��v���~��
����:���7���N�P�W�s�N��8�y��N���i]��!2��P   P   ܃�7�R��$1�\� �ށ �*k0�z�Q�d��!{��.�ٽ��
��U*��mF��iW�P�W�"�F���*�{'�n�ڽ����P   P   �v����e�,�<�N %�5�_�$���;�GOd��d��U���T,�����0��mF���N�N�F��X1�D��Ѱغ�P   P   ����6Nu���F��v)���u����(�ŊE�Hs�̱��@7ýJK�����U*���7���7���*���h���T�ĽP   P   �r����}��JN�Ow-�zC�������L,�2�L���{����@7ýT,��
��:�9����n#���ĽP   P   c��� ~���P���/��N�,���P��s��X.�
�N���{�̱��U���/�ٽ���.�`V�A�����ڽ���P   P   )�����u���N���/�!W�ɟ�k2	�y"�Q��X.�2�L�Hs��d��!{���~��zBν�2Խ�νEs��Ъ��P   P   ���9bf�AqG�f�-��������R��y"��s��L,�ŊE�HOd�e���v��Ԡ�Yy��w����n��|[��P   P   m�i�*8S��O=�t*����l�c�	��R�k2	��P�����(���;�{�Q���g���{����׸���[���3}�P   P   �K�?���1���%�������l����ȟ�,�����u��_�$�*k0�j�=�x�J�� U�Y[��S[��U�P   P   ߜ1��J,�_�&�X�!��)����������!W��N�yC���5�ށ �m�%��F+���0�,�4�ڀ6�^5�P   P   ��Z��V@�x��X�!���%�s*�f�-���/���/�Nw-��v)�N %�\� ����T����]�R���
�P   P   ���w��	��V@�^�&���1��O=�@qG���N���P��JN���F�+�<��$1�G�%�0��P�Pg�����P   P   ��6��w��Y���J,�?�)8S�7bf���u�� ~���}�5Nu���e�7�R�v�>���+����p�n��l�P   P   냹������ռ�Q���V�h�5� \��2������ك���1���f���L���u[��<5�8��W�����Լf]��P   P   e]���`��9�Ҽ����4�Z�B��v��P���յ��νu�ܽ�ܽ�qνS���i&��#�u�f�B�i������ҼP   P   ��Լ ɼ1�Լ����(���J����8����ս4��������)�W����ս�|��(���J�:������P   P   W���:�ڼ�ڼ-J��ŵ�%�I��H���˴�R���v�"�-��@=��B=�T�-�\��
�W�������J�i�P   P   8��O�������
���q���A�����~������n��E�.c���n�4Qc���E���Sm��W��(��f�B�P   P   �<5�������)#���n�LU4�xt������뽞(��mN��ez������
��t�z���N���
콙|��#�u�P   P   �u[���$��������e���#��Y�)����ӽ�����D��z��z��Z���t���u�z���E�]���սi&��P   P   �h>���h� �gR ������<��ր��(���
���,��;b�M���QК�Z����
��4Qc�T�-�X���T���P   P   �L��AqW�j�"�����n���#��!�(JU��֒���̽o����;��{m�M����z��������n��B=�)��qνP   P   �f��Σk��70�J��.������Ϯ
��[.��h�-����ڽ�v���;��;b��z��ez�.c��@=�����ܽP   P   �1��\w�Յ9�1����<伛<�9j�K7�	t�-=���ڽp���,���D��mN���E�#�-���w�ܽP   P   ۃ��(2w�b =���o�󼩥ڼ��ټ����9���:�	t�-�����̽�
������(��n� w�6����νP   P   ����!l��9�M$���� {ּAR̼�ռ���9�K7��h��֒��(����ӽ�뽐��T�뽬ս�յ�P   P   �2��C�W��0��U�	�����ּ�Aȼ�Ǽ�ռ���9j��[.�)JU��ր�*������ ~���˴�:����P��P   P   \�!?���#��y�8����ۼt=ͼ�AȼAR̼��ټ�<�Ϯ
��!���<��Y�xt������H������v�P   P   j�5�{�%�dR�������aE漨�ۼ��ּ�zּ��ڼ<伖��#������#�NU4���A�'�I��J�\�B�P   P   �V�֙�ߺ������������7��������n����.����n��hR ��e��n��q�ǵ�*���4�P   P   �Q��F������b���������y��U�K$���0��I�����h� ����*#���
��/J���������P   P   �ռT�ۼ	;����޺�cR���#��0��9�a =�ԅ9��70�j�"��������������ڼ2�Լ;�ҼP   P   ����O�ɼT�ۼE���ՙ�z�%� ?�A�W�l�%2w�Zw�̣k�?qW��h>���$���P���;�ڼ ɼ�`��P   P   Q>�`�M��i|�"g��4��8p�lH��}|����9:��������US����{�=�G�������8쥼L�{��rM�P   P   �rM��5M��<w�Ѳ�������(��j�1���25Ľ%.�,���ͯ��� 罎�ý�y��۷i�}�(����k���m,w�P   P   K�{��`��1{��C��_"�j/2�F���Z�������a��t-��76�k-�Y�w�𽭄����� k2�k��k���P   P   8쥼� ��׃�:G����켁�1��*��m�½k����5���_�
3z�x;z��`�6�B	�Lý<���!k2����P   P   ����裼���1����߼$�'�f��[½�����H�{<��@���w1��Q��o���lI�Sa�Lý���}�(�P   P   ����мV������ڌμ���^�g��[��$S���H�����[���iϾ��Ͼ�����n���lI�C	�����۷i�P   P   =�G����dQ��83��]���i���E�1����{�4�T�������޾���M߾�����o��6�x��y��P   P   ��{��e#��N߼�a��Ō���ݼ�i!�L�x�����l��S@^����ξ_�����ϾQ��`�Y���ýP   P   VS����B�l��㼼����<��o  �	@��X���A佁�+�Ax�8 ���ξ��޾�iϾx1��y;z�k-�� �P   P   ���<�\�
&���˼=Ϣ��䡼�:ɼ���3?Y�u����z���D4�Bx�����[��@���3z��76�ϯ��P   P   ���5�k������ؼQ����+��b���Gռx��P�g�?���z����+�T@^�U�������|<����_��t-�.���P   P   ::��'�k�"M"������M���q��Ed��>�ܼT*�P�g�u����A�l��|�4���H���H���5��a�'.�P   P   ���&]�R$��0�c��t���fo����
��>�ܼx��4?Y��X��������%S����m�����45ĽP   P   �}|��iC����
�ټ~���@���n|f�8We����Ed��Gռ���	@�N�x�2���[��[½o�½\���3���P   P   lH�}$�e|��~ͼ�7��f�����q�m|f��fo��q��b����:ɼp  ��i!���E�a�g�f���*��G��� j�P   P   ;p��f���ᾼu񤼱s��f���?���s���M���+���䡼�<���ݼ�i����&�'���1�l/2���(�P   P   7��YPѼ<��Ó���D��t񤼇7��|���a����P���=Ϣ����ƌ��_��܌μ��߼���c"���P   P   $g��%���.��y��Ó���ᾼ�~ͼ�ټ�0�����ؼ��˼㼼�a��93�����1��=G���C��Ӳ��P   P   �i|��Ȅ��x���.��;���d|����P$� M"����	&�k���N߼dQ��V������׃��1{��<w�P   P   a�M��a��Ȅ�$��WPѼ�f�z$��iC�&]�$�k�2�k�:�\���B��e#�����м�裼� ���`��5M�P   P   f��:Tp�9��,�����4����",�]\m����T��@����笽ྕ�U�l��+���⼈��� ��T*���9P   P   ��9���96��Eh�����A���V�Ą��Usҽ�5�T��u��w�V5ҽ>P�� �U����������X��P   P   �T*��C�՛(�N~�♼�'� �t��r�����>%3��U��:c�#�U��3����Y���'�t�u��������P   P    ���`��^�sC�Ρ����R>�/�н��~�b�䒾�򨾲���T�����b���G1ѽ���v������P   P   ����I���Ѣ�t����ー)���s��н�D(��M��kG���R徭�����1���������(�H1ѽ'�t����P   P   ��⼳"b����[����{^�'�߼�S�c껽������k�¾R��]�$�h�$��M���þ���� ��Z����U�P   P   �+�Fc���`9�}S�516�DG��B�(��o�����a�N\��܍��6�M��H7��M�1�����b����?P��P   P   W�l��4��󶃼�Q�6Q����=����h��_Ͻ�	1�z�����㾜�#�Z�L�M�h�$���U����3�X5ҽP   P   ᾕ�B�%� |���[:�>���`6����� "�X��ec����R��$��~�����#��6�^�$���������%�U�x�P   P   �笽V)F��Tּb_�X������sX�H�мo�A�{���d�0`��$�����܍�S���R徾��:c�v��P   P   B����X�J�����!��G�����hw�\�켋�S�}��d���R�{���O\��l�¾lG��䒾�U�U��P   P   V�� Y�?9������
��`��ץ�����;{��������S�{���fc���	1�
a�����M����b�@%3��5�P   P   ���1�F��:�����k��R.�[U���K�;{��]��p�A�Y���_Ͻ�������D(������XsҽP   P   a\m��?&���׼]��)����h�����[U������hw�I�м� "���h��o��e껽�н1�н�r��Ǆ��P   P   &,�A������g1b�%M����;9�f��P.�ץ����sX�����=��D�(��S��s�V>��t��V�P   P   ��=ó��o����>�����bĻ������h���`���G�������`6���GG��+�߼+�����'�D��P   P   �4����d�+�<����"[����#M�&����
��!�W��?��8Q�916��{^��ーҡ��
♼����P   P   �����������	������>�b1b�Z���������__��[:��Q�~S�a���}���xC�T~�Jh�P   P   �,�Mf�z�������'�<��o�������׼�:��;9��G���Tּ�{��󶃼�`9������Ѣ��^��(�B��P   P   1p�9![R�Mf������d�9ó�<����?&�.�F��Y��X�S)F�A�%��4��Ec���"b�	I����`� �C�U��9P   P   ��<.a}<&I<��;8�����
���S��揽�Ҭ�����������\R��������4���;�.I<|�}<P   P   |�}< �}<MCM<=��;� ��� ���e6�0ɗ�}�۽�]�ȿ �� ��=���۽ꘗ�;6�V/���X�����;	vL<P   P   �.I<�(i<l$J<��;�Y���ɼ0[�������RQ��e��&B��b��dKQ����(��,�[�H�ʼwN�����;P   P   ��;9�;<��<<�0�;)o���sȼ�Gh�\�ٽ�6��؊�9 �������ᾞE��
��%s6��NڽO�i�H�ʼ�X��P   P   ��4�'1�;��!<�U�;�#�;�{tY��ؽ�B�j8�������'���;�b'��R��	ԡ�2C��Nڽ-�[�W/��P   P   ���o��8��;�b�;e�9� x�3^3���q�4�a����,�BiS�ډ�	��RT����
ԡ�%s6��(��;6�P   P   �����t6;+*�;lnE;s
��� ��0���K��������8�R��|�������RT��R��
����똗�P   P   �\R�-����,�~�;��;cs�
�����M���׽�ZN��黾�s%��刿U躿|���	��b'��E��eKQ���۽P   P   �������\�3D ;QF�;L�2;������S��v�
���~���޾H�9��刿�ډ���;����b���=�P   P   �����$���k�H��x�;�c�;�~/9	n^��R�������������޾�s%�9�R�DiS��'����'B��
� �P   P   ����Y;���L2�V�;E�<�c�;�Y
�����M95�,�������~��黾����,�����; ���e��ʿ �P   P   �Ҭ�b�;�����wӈ����;��<,�<�ʬ;�Lb�9ۛ�N95����w�
��ZN�����b���k8���؊��RQ��]�P   P   �揽�#%�R���������;&�<�D0<[�<�K�;�Lb������R�S����׽�K�s�4��B�6�����۽P   P   S�.:��,<n���:�3H�;��<�"7<E�8<[�<�ʬ;�Y
�n^���󼨧M��0�� ���ؽ`�ٽ���3ɗ�P   P   ��@�������5��/R�;�<M�-<�"7<�D0<+�<�c�;,~/9�������� �7^3�tY��Gh�0[��e6�P   P   ���f����9�l�;���;�&�;�<��<'�<��<E�<�c�;@�2;vs�!s
�� x�A�tȼ�ɼ� ��P   P   :8�;�29);A��;��;���;4R�;9H�;���;��;X�;�x�;NF�;��;ZnE;��9�#�:o���Y��� ��P   P   ��;��;l�;��;E��;z�;�4��y�:����mӈ��K2���6D ;}�;'*�;�b�;�U�;�0�;��;2��;P   P   &I<��:<�S<�l�;B9);��9����#<n�N�����������k�Y��,��t6;��;��!<��<<i$J<ICM<P   P   -a}<5�h<��:<��;*;�]��:���':���#%�_�;��Y;���$�����+�������8&1�;8�;<�(i<��}<P   P   ^=�=z�<H��<8�W<��g��枼�\(�񬀽����ꄯ�����@[����'�� ����W��-X<֞�<sR�<G�=P   P   G�=�=Hx�<���<.4<�����:R���)ڽ�F�5.+�"+�J#��ٽ&������.�2<��<�<P   P   sR�<��<M��<�)�<�''<!�-�x�0��������`�h�i���Nܡ�ɟ��8�h����ֹ�NZ1���0�-f$<��<P   P   ֞�<zF�<���<��<37<`j+�u�?�V�ֽ��E��2�����3�����N�辖{���-F�5�׽qCA���0�.�2<P   P   �-X<Ꮏ<�k�<���<�7]<�ػA�.���ս��T� ¿�D�Wi�	R����i�V��\����&V�5�׽NZ1����P   P   ��W��:�<%��<�{�<'ӆ<EϚ�^��,Q���7D�����2�:��{h޿H�޿�!��5N4�\����-F�ֹ��P   P   � ���-�;$5�<ϲ�<_6�<;��;�і�GJ�����*������+|�������+�h�	��!��V���{�����&��P   P   ��'��D��7�S<���<���<�|[<M����F"�-eս�d�1v�vf� ܿ� +���+�I�޿��i�O��:�h��ٽP   P   A[��VR��ܟ�;�=�<�Ȱ<��<K��;h�����x����.둾����U�� ܿ���}h޿
R�����˟��L#�P   P   ����o�*Ĺ�\p<�{�<��<0�x<��:��޼�����I'�Iʞ����vf�,|��:��Wi�5��Oܡ�"+�P   P   섯����#$��X�@<hϥ<�.�<q�<%L<kv������*���I'�.둾2v御����2�D����k���7.+�P   P   ���������߻��$<�9�<�~�<a��<�͡<��1<�ݷ������������d�+�����¿��2��c�h��F�P   P   ����j������S'$<#��<�ؿ<o��<��<��<��1<ov����޼��x�/eս����7D���T���E�����)ڽP   P   �\(�����s��H?<�k�<P�<��<���<��<�͡<#L<m�:l����F"�IJ��/Q����սZ�ֽ����>R��P   P   �枼�C��j�;�tm<r?�<���<���<��<o��<a��<q�<-�x<@��;^����і�b��F�.�z�?�~�0���P   P   \�g�f�;�;Q<�c�<�S�<��<���<P�<�ؿ<�~�<�.�<��<��<�|[<+��;�К�"�ػnj+�0�-���P   P   0�W<聃<X��<p�<Bޭ<�S�<s?�<�k�<%��<�9�<iϥ<�{�<�Ȱ<���<\6�<$ӆ<�7]<)7<�''<.4<P   P   E��<�<�Y�<A}�<p�<�c�<�tm<�H?<Y'$<��$<[�@<�\p<�=�<���<Ͳ�<�{�<���<��<�)�<���<P   P   z�<���<]�<�Y�<Z��<<Q<z�;ds�������߻$��r)Ĺ��;8�S<$5�<$��<�k�<���<K��<Fx�<P   P   �=���<���<�<끃<x�;wC������b�뼤�����j�SR���D���-�;�:�<���<yF�<��<�=P   P   F�Q=��M=F�@=��'=�d�<�)�<�TS�D�ټ��M��;��MI������7M�1�ؼ��L��]�<G6�<(}'=s{@=پM=P   P   پM=9�M=q�A=�^&="i�<�%<����B^��ȽЉ���)�	{)� b��ǽ��]�A���
�#<�|�<W�%=�yA=P   P   s{@=`�H=b�@=Z�&=G�<��;/�%����	���n�������j��n���{ڣ�b����;���<W�%=P   P   )}'=gc==�==�C(=���<���;�M�p�ý>�F������ �#�"��"�(� ��򫾞vG��Ľf���;�|�<P   P   G6�<s)=�86=/(*=�x =5P,<��⼼�½4,X���Ͼ��7�����Η��g]����8�+�о�Y��Ľc��	�#<P   P   �]�<O�
= �(=gg)=#=�+�<^�������>E�cϾ< Q���ÿ"���A��1ſ��R�+�о�vG�{ڣ�B���P   P   ��L����<�=��$=��=0e�<A�:�W�a�������96�}�¿uN<�1r�P�=��1ſ��8�������]�P   P   5�ؼuh2<=�<��=�Y=�F�<�A<ϼ̼��½�xj�s���"������q�2r��A�h]��(� �
�n�
�ǽP   P   �7M�(#�]ӷ<K�=�[=�=�̽<?����D��
��ș�����������vN<�#��З���"�k�"b�P   P   ����g�� |<���<}!=��=�a�<�H�<�M�b����&%�騾���#���¿��ÿ����%�"� ���{)�P   P   PI��w��H'<�F�<f�=V=$%=�/�<Ph:<�ٜ�i}���&%��ș�u����96�> Q���7��� ������)�P   P   �;��[`��n�<8;�<nE=��=��=�4=���<�,<�ٜ�c����
��xj�����fϾ��Ͼ�����n�҉�P   P   ��M�_�i�=�%<���<�)	=��=�	=�=k=���<Mh:< �M���D���½c���>E�7,X�B�F��	��ȽP   P   O�ټ/�+�hz<%��<B�
=�w=z�=^�=�=�4=�/�<�H�<�?��ּ̼@�W������½t�ý)���B^�P   P   �TS�j_0<~��<��<.=�B=s[=z�=�	=��=$%=�a�<�̽<wA<:A�g�����⼧M�:缲���P   P   �)�<���<(�<��=i=�=�B=�w=��=��=V=��=�=�F�<,e�<�+�<'P,<���;Ş�;�%<P   P   �d�<��
=rD=��=�=i=.=B�
=�)	=nE=f�=}!=�[=�Y=��=#=�x =���<�F�<i�<P   P   ��'=^[)=Cw(=ԉ#=��=��=��<'��<���<:;�<�F�<���<J�=��=��$=fg)=-(*=�C(=X�&=�^&=P   P   F�@=�W==��5=Cw(=sD=+�<���<'hz<F�%<v�<N'<� |<^ӷ<=�<�= �(=�86=�==a�@=q�A=P   P   ��M=�H=�W==_[)=�
=���<u_0<��+�P�i�T`��q���g��'#�xh2<���<O�
=s)=gc==`�H=9�M=P   P   �t�=<��=�Z�=�{t=��K=�?=�s<�F���
��5X�<�u���W�x�	����t<�==�K=t=�(�=I��=P   P   I��=ɖ�=�ӆ=�zs=LD=���<�V\:�j��>��A' ��]�!����ȧ����2�a:���<�pC=��r=��=P   P   �(�=��=�\�=A�s=(A=eb�<�N"�������c�F���\ʧ��藾u�b�ej�����pk$����<�@=��r=P   P   t=�b�=x��=w�t=`�D=1��<�b��T��\�9�3ʦ�:���� �p� �9'��	����9������h����<�pC=P   P   �K=��t=0��=��u=�#M=6/�<���W�� VK��˾�5�K����{��P݊���6�Ĥ̾�L����qk$����<P   P   �==f�U=9�r=�Ms=r�V=��=�i�:.~�1�7���ʾmO�l����O���� ¿�P�Ĥ̾��9������a:P   P   �t<B*=3�\=�l=U^=|�,=�"�<��l��<ˤ�YE4��d���[7��0k� �8�� ¿��6�
��ej����P   P   ��9-�< X@=�__=�`=]oB=���<s�������|�^�������B��V�i��0k���Q݊�:'��w�b��ȧ�P   P   z�	�\�l<`�=,N=�+\=��O=L�"=�Ӏ<�������˔����Ϙ��C���[7��O��{��r� ��藾#���P   P   ��W�k�;�� =��;=?�S=�T=��==�=�;�%M����2��������d��n���L���� �^ʧ�^�P   P   A�u�^��q��</�+=��I=!S=aeK=9�.=c��<r'G�*�i����˔�����ZE4�oO��5�=���H����P   P   �5X�⊢�K��<��!=� B=�#O=g�O=OD=�t%=ǈ�<|'G��%M�����~�^�>ˤ���ʾ�˾5ʦ��c�C' �P   P   ��
�?�;�9�<l�!=?=�:L=P=�HM=_IA=�t%=b��<ָ;������o��4�7�VK�`�9����>��P   P   �F���j<�Y =^@+=��A=|L=1�O=��O=�HM=ND=8�.=
�=�Ӏ<������.~��W���T�����k�P   P   �s<R[�<O=�!;=JhI=��N=uO=1�O=P=f�O=aeK=��==K�"=���<�"�<Yi�:+����b��N"�aU\:P   P   �?=N*=S�?=��M=��R=��Q=��N=|L=�:L=�#O=!S=�T=��O=[oB=y�,=��=./�<*��<]b�<���<P   P   ��K=�oU=��\=O�^=*	[=��R=JhI=��A=?=� B=��I=>�S=�+\=�`=T^=p�V=�#M=]�D=%A=JD=P   P   �{t=��t= �r=�Kk=O�^=��M=�!;=_@+=l�!=��!=/�+=��;=,N=�__=�l=�Ms=��u=u�t=@�s=�zs=P   P   �Z�=�x�=�x�=!�r=��\=T�?=O=�Y =�9�<N��<s��<�� =`�= X@=2�\=8�r=0��=w��=�\�=�ӆ=P   P   <��=��=�x�=��t=�oU=P*=X[�<��j<w�;Ɋ���]����;_�l<:-�<B*=e�U=��t=�b�=��=ɖ�=P   P   �=L�=k3�=��=�u�=qqY=a�=���;i
�����b+9��.����X�;�=�nY=�:�=�8�=��=o�=P   P   o�=/	�=���=�j�=�P�=�3C=o�<����𶈽���1������:⽺އ�����B�<8�B=���=��=iy�=P   P   ��=�w�=�,�=k~�=B�=��5=�O<�J?����T�Ц���Ҟ�J|����S�����]u>��<-�4==��=��=P   P   �8�=�ƨ=���=鯟=a��=b(6=[q�;XՀ���*��ܝ����,��}�ɝ�)w*�P�����;-�4=���=P   P   �:�=��=5�=��=?��=��D=�<����O<�����6 &�Rns�����c�s�cd&�M4����<�Q����<9�B=P   P   �nY=5��=!�=�^�=vK�=^�[=v��<�t:�)�;
���:�ف��K�߿~�S��n�;�N4��*w*�^u>��B�<P   P   �=�p=��=��=*��=�{r=��=<=�����8$��)�$��͟�:_���'�bX�S��dd&��ɝ��������P   P   �X�;�8=2,�=kM�=͞�=�9�=m�;=��<#���	&P�4����p���ݿ�,'���'��e�s���S��އ�P   P   �����<͙\=l��=ϓ�==S�=�_=�� ={���.$ܽ��=�B̉���ݿ;_�M�߿����.��L|���:�P   P   �.�[�<z�:=pp=���=G�=��r=R�>=؛<_���	��ӛ��=���p��͟�ځ��Uns�����Ҟ����P   P   g+9�j� <j�!=h8]=p�v=P�}=�x=�4`=Ź&=.C><'2.���	��5��+�$��:�8 &���Ҧ��3��P   P   ����<��=
R=��k=�t=H]u=ҝm=��U=d�=+C><
_�1$ܽ&P�9$��=
�������ܝ�T����P   P   t
��k��<i�!=r�Q=I]g=��n=��p=�p={�i=��U=Ĺ&=؛<����&������)��O<���*�$�������P   P   x��;0��<�5:=��\=�sk=n�n=K�n=6o=�p=ҝm=�4`=P�>=�� =�<H=���t:����]Հ��J?�����P   P   ^�=O�7=Q\=�p=�9v=�$t=c\p=K�n=��p=G]u=�x=�r=�_=j�;=��=l��<�<(q�;�O<o�<P   P   nqY=$p=��=�\�=?3�=�|=�$t=m�n=��n=
�t=O�}=F�=<S�=�9�=�{r=[�[=��D=^(6=��5=�3C=P   P   �u�=r��=�ޏ=��=��=?3�=�9v=�sk=I]g=��k=n�v=���=Γ�=̞�=)��=uK�=>��=`��=A�=�P�=P   P   ��=8��=��=<��=��=�\�=�p=��\=r�Q=
R=g8]=pp=k��=jM�=��=�^�=��=诟=j~�=�j�=P   P   k3�=[�=�4�=��=�ޏ=��=Q\=�5:=j�!=��=j�!=z�:=̙\=2,�=��=!�=5�=���=�,�=���=P   P   L�=}��=[�=9��=r��=&p=Q�7=5��<q��<�<q� <]�<���<�8=�p=5��=��=�ƨ=�w�=/	�=P   P   :}�=<��=?W�=ҭ�=Vd�=�-�=�==�S�<�;�y������b���B��V.�<rG>=6�=%�=�Q�=G�=���=P   P   ���=���=�J�=�y�={��=*f�=��=A�%���{��#�#k�x%�h�ཱི�x��g�k�=Rc�=5�=K�=L��=P   P   G�=\/�=(K�=C��=�֩=N_x=�<��������]����Wh������\�U���g����<Dx=�[�=K�=P   P   �Q�=@�=xL�=R��=�Ϊ=�y=ʱ�<�If���/�Q�����>������Y���ݦ���.��Nd�!�<Dx= 5�=P   P    %�=B�=�\�=���= �=�5�=���<o�d���C�2;��,�Xq���|$q�/�,�\�̾�C��Nd���<Sc�=P   P   6�=o$�=Dp�=İ�=|�=�F�=K.
=-��An.���̾wB@�����Xǿ�ǿ�����K@�]�̾��.�g��k�=P   P   sG>=I��=H$�=l@�=[��=��=i�A=��O���+��<#,��=���`� V�������0�,��ݦ�W����g�P   P   V.�<�l=�=GV�=W��=�ə=��o=�ŧ<.Xr��]Z�����L�o��&ƿT�V��ǿ~$q��Y����\���x�P   P   G���*=�A�=��=l�=җ=�ǅ=�R/=�\軆�۽�Օ��I�h����&ƿ�`�Yǿ�󇿋�����j��P   P   h����J�<K�a=z�=rr�=�Ր=C��=<�e=hz�<����������I�M�o��=������Xq�@��Xh��z%�P   P   ����2�<58E=�|x=�c�=î�=��=�{=FJ=.Z�<������Օ�����>#,�yB@���,������%k�P   P   �������<��:=�j=��z=��~=�k=�|=�$n=�?=,Z�<��載�۽�]Z�+����̾2;T�����]��#�P   P   �;��<��D=��j={Uu=ku=�!t=v=��w=�$n=EJ=cz�<�\�5Xr�U���Dn.���C���/������{�P   P   �S�<��)=*Ya=T_x=��z=n�t=�o=Q p=v=�|=�{=9�e=�R/=�ŧ<	��6��z�d��If����^�%�P   P   �==�l=�)�=�Y�=�8�=�K~=��s=�o=�!t=�k=��=B��=�ǅ=��o=d�A=F.
=���<���<�<��=P   P   �-�=���=���=�=0�=�G�=�K~=m�t=ju=��~=®�=�Ր=җ=�ə=��=�F�=�5�=�y=J_x=(f�=P   P   Ud�=�O�=1�=�3�=&��=0�=�8�=��z=zUu=��z=�c�=qr�=j�=U��=Z��={�=�=�Ϊ=�֩=z��=P   P   ѭ�=���=��= �=�3�=�=�Y�=S_x=��j=�j=�|x=z�=��=FV�=k@�=ð�=���=Q��=B��=�y�=P   P   ?W�=La�=
v�=��=1�=���=�)�=+Ya=��D=��:=48E=J�a=�A�=�=G$�=Cp�=�\�=xL�='K�=�J�=P   P   <��=�`�=Ma�=���=�O�=���=�l=��)=�<���<�2�<�J�<�*=�l=H��=n$�=B�=@�=\/�=���=P   P   ���=l��=�H�=�V�=�y�=Ρ=�B\= ��<r�@�2Q��/E���a~6�#�<U�]=��=�3�=
��=��=���=P   P   ���=���=���=�;�=���=ߙ=>�#=1�6��
��2;�&f3�W�2�4	
�Xo����&��%=��=mD�=��=�.�=P   P   ��=���=f5�=lD�=,C�=���=r��<�\8�_[��A��];þ_-پ�b¾�
��UA�3�,@�<\	�=	��=��=P   P   ��=9��=��=�e�=E��=K�=��<	爽��[�Q�ؾ��'�׶Q��MQ��&���־�UY��M���7�<\	�=mD�=P   P   �3�=/C�=I��=���=���=���=�(�<C����Dv��`���j�����Ժ�����r�i�KT��t��M��,@�<��=P   P   ��=��=���=��=Zc�=��=�<'=KY3�bwZ��������2ӿ�A�/�w~ҿ�悿KT��UY�3��%=P   P   V�]=ئ=���=���=3V�=���=Pi`=֓��	��4׾}:j�(�ҿ�{�7�.��P�w~ҿs�i���־UA���&�P   P   $�<*��=H�=�w�=/ٯ=��=�3�=X��<_��_���&��������.�7�.�0������&��
��Yo��P   P   c~6�ҳ9=��=�l�=�2�=�3�=M/�=-R>=�n�/������P�$k�����{��A��Ժ��MQ��b¾5	
�P   P   ��1P�<h=(̇=��=H�=���=bl=�[�<�6�O0�e=׾��P����)�ҿ�2ӿ���ٶQ�b-پZ�2�P   P   �/E��n�<E�E=X�o=q�x=�y=�,z=��r=oJ=�Ҧ<�3;�O0�����&�:j�������j���'�_;þ)f3�P   P   7Q��՗<3�8=��]=s�a=�^=�^=%�c=#a=�>=�Ҧ<�6�1�a���4׾���`�U�ؾ�A��5;�P   P   ��@�}�<�EE=Д]=PyY=�uN=�I=j�O=��[=#a=	oJ=�[�<�n�c���	�gwZ��Dv���[�d[��
��P   P   ���<D�8=��g=��o=Ŗa=rNN=ݮA=yB=i�O=#�c=��r=_l=)R>=L��<���VY3�J���爽�\8�R�6�P   P   �B\=n>�=ܐ�=���=k_x=1�]=I=ܮA=�I=�^=�,z=���=K/�=�3�=Ki`=�<'=�(�<��<d��<8�#=P   P   Ρ=Ӧ=��=]�=��=~�x=1�]=qNN=�uN=�^=�y=H�=�3�=��=���=��=���=K�=���=ߙ=P   P   �y�=���=��= q�=V�=��=j_x=Öa=NyY=p�a=m�x=��=�2�=-ٯ=1V�=Xc�=���=C��=+C�=���=P   P   �V�=��=��=���= q�=]�=���=��o=Δ]=��]=T�o=&̇=�l�=�w�=���=��=���=�e�=kD�=�;�=P   P   �H�=m�=k�=��=��=��=ܐ�=��g=�EE=1�8=C�E=h=��=F�=���=���=H��=��=e5�=���=P   P   l��=��=m�=��=���=Ӧ=o>�=F�8=}�<�՗<�n�</P�<ϳ9=)��=ئ=��=.C�=8��=���=���=P   P   թ >���=��=aL�='��=Υ�=��Z=C~n<��߼`�y�����w�}ؼ�6{<e�\=�ժ=�b�=���=�	�=hU�=P   P   hU�=C�=�m�=��=��=p|�=q� =!�ü��׽��@���w���v���>�?�ӽ�뷼5�#=�֥=�_�=��=���=P   P   �	�=���=�f�=��=#t�=���=t�<o|��"S��xþ1�
����7
�n��w�O�zW����<n�=~
�=��=P   P   ���=���=��=�P�=���=��=,�<���
�������z�D����V��iy��$�$͕�����,�<n�=�_�=P   P   �b�=l[�=��=��=��=dX�=�:�<�´Ӫ�sTE�;,��#�J�����"���<=C�{���������<�֥=P   P   �ժ=��=\<�=݊�=�G�=�̫=��$=噄�Y$����D��9Ϳk�*�V�\��-\�տ)���˿<=C�$͕�zW��6�#=P   P   h�\=@©=n��=��=f^�=��=�;_=z޴��VP�A������>b*��u{��H����z�ֿ)�"����$�x�O��뷼P   P   �6{<��}=l=�ܦ=?�=��=���=f��<[ҽ�K��Koy�����m\�W���H���-\����ky�n��@�ӽP   P   }ؼ�=��|=�#�=��=��=1�=؉$=��˼6�<�3�	�t
��	���m\��u{�X�\�L���V���7
���>�P   P   �w��-�<i@=�\=W�^=u�_=x_=fD=���<B#n�2�s����t
�����?b*�m�*�$�G�������v�P   P   ���O�;\Q=L�0=�,=�(=�K.=w4=�=-x<����3�s�4�	�Noy������9Ϳ>,����z�4�
���w�P   P   f�y�y�;Wr=�(=�w
=ض�<V"�<Y�=� =� 
='x<F#n�8�<��K��C����D�wTE�����xþ��@�P   P   ��߼��<K=�=Z7�<��<A'�<k�<e� =� = �=x��<��˼`ҽ�VP�\$���Ӫ��
��"S���׽P   P   /~n<�x=�?=�0=�Q
=�r�<�'�<�)�<h�<V�=s4=fD=҉$=W��<�޴�완��´��v|��5�üP   P   ��Z=##}=�u|=��\=Ah,=��<Z�<�'�<<'�<N"�<�K.=x_=+�=���=�;_=��$=�:�<�+�<t�<k� =P   P   ͥ�=!��=�؞=�"�=f�^=׹'=}��<�r�<��<ζ�<�(=o�_= ��=��=��=�̫=bX�=��=��=n|�=P   P   &��=���=J�=��=W׋=e�^=@h,=�Q
=S7�<�w
= �,=P�^=��=?�=c^�=�G�=��=���="t�=
��=P   P   `L�=L��==��=u��=��=�"�=��\=�0=�=�(=G�0=�\=�#�=�ܦ=��=ڊ�=��=�P�=��=��=P   P   ��=�=�s�==��=J�=�؞=�u|=�?=I=Tr=WQ=d@=��|=j=k��=Z<�=��=��=�f�=�m�=P   P   ���=>��=�=L��=���=!��=$#}=�x=��<y�;O�;�-�<�=��}=>©=��=k[�=���=���=B�=P   P   �>�
>�p >I�=��=���=Y�8=��к�X�ɠ��6��;����S���%���:=�Ϥ=D�=R��=[" >��>P   P   ��>t�>{>��=���=�)�=�:=ٙ3�A�O?��ܞ��b��w������,�H�=���=;%�=(p�=��>P   P   \" >,2>-Y >��=���=;̢=�|�<j����/��"���I>�b�V�U.=�# ��ۉ�o���ߠ<�4�=���=)p�=P   P   S��=��=��=G�=w��=��=�9P<�=��ʾGV�g���!�{�俜��D�S�y�ƾ�6 ��}`<�4�=<%�=P   P   D�=|a�=M+�=��=��=��=��<��0侌M����b�@��J[�E�?����#���E���6 ��ߠ<���=P   P   �Ϥ=��=�>�=���=¸�=�ӥ=��=�{���ȾO��n��+�z�ʇ��AK��ֻy����#���y�ƾo��K�=P   P   ��:=蕙=�=���=��=��=hk==[�*��k����T��C��z��������C��ֻy����E�S��ۉ��,�P   P   ��%��SI=�)�=Mi�=�ӄ=�o�=qM=���9X���%�SU���)@�Xs���������BK��F�?����$ ����P   P   ��S�!��<�|)=|,4=;q2=T6=",-=�j�<��L��}��}<�u�*[�Xs�����ˇ���J[�}��W.=�x��P   P   <��呻=��<�}�<�>�<TR�<?l�<z��<W1�麽Y4���/U�v俵)@��z�.�z�e�@��!�e�V�e��P   P   8�⽬���G�<�:<�Va;��9:�;�$<��<�F��$ܽZ4���}<�UU���C�q����!g���I>�ߞ��P   P   ̠�����V�?;��6:h/�oǄ�����*�
�ʔ�:�
�;�F��麽 �}��%���T�Q���M��GV�%��R?��P   P   ��X�Ꝼ�a<��3:��]���мV��V�ͼہR����:��<�1���L�[���k���Ⱦ6侣ʾ�/��A�P   P   t�к�˧<ò<¢<��BѼ�!�ٛ�[�ͼ9�
�Ѯ$<m��<�j�<��9h�*��{�����=�r����3�P   P   V�8=cnH=U7)=�F�<��[;�"�������!�^������|;/l�<,-=iM=`k==}�=��<�9P<�|�<�:=P   P   ���=U��=H�=3>4=�K�<���9�"��IѼ �м~Ǆ���9:BR�<K6=�o�=��=�ӥ=��=��=9̢=�)�=P   P   ��=!A�=T�= w�=0�1=�K�<��[;���]��/��Ua;�>�<1q2=�ӄ=��=���=��=u��=���=���=P   P   I�=���=���=J��= w�=2>4=�F�<��<8�3:��6:�:<}�<r,4=Ii�=���=���=��= G�=��=��=P   P   �p >�==��=���=T�=H�=S7)=ò<ta<��?;(�<+��<�|)=�)�=�=�>�=K+�=߿�=-Y >{>P   P   �
>Le>�=���=!A�=U��=dnH=�˧<	Ꝼ�������9呻��<�SI=啙=��=za�=��=,2>t�>P   P   ��>1}>f��=+��=�%�=z�=Hl�<��ɼm��������������g���Z��<f(�=��=m��=� �=�I>P   P   �I>�h>�C >���=��=��=Ʃ�<�����E8��d�ƾ��ž-0��V5� �|���<ݙ=Iq�=f��=���=P   P   � �= ��=<��=���=���=�$�=_L*<Ҍ�\S��Q����c����I�b����˥��o�7><Y��=�,�=f��=P   P   n��=���=�=�=~�=�:�=��=��;���<���@��C�׿b���h��	ֿ�o}��.꾤+����;Z��=Jq�=P   P   ��=�]�=z��=� �=S��=�~�=�]6<+��*t�G����}���l�u߆���k��?�'�������+�>><ݙ=P   P   j(�=��=h�=�a�=��=gb�=���<ތ����>����5�/ܙ�х��U��=���s4�(����.� o���<P   P   j��<:d=Iv=�v=e�w=�Vg=x�<0H{�P8��	�~� ��%���������������=���?��o}�̥����|�P   P   Y���۷�<��=`��<�
=O�=M��<a#���04�F��u@ֿal��h����������U����k��	ֿ���V5�P   P   �����l6��I;���9��]8�:��;���Bg��Q֘���a��窆��h������Ӆ��w߆��h�L�b�.0��P   P   ���W+�+z��o2�w3�2�����%���F�"�����þJ���bl�'���0ܙ���l�d�������žP   P   ��8wv�}�*��$P�����:y�������jK�>d#��&l�
��þ��a�w@ֿ"����5��}�G�׿��c�g�ƾP   P   ���� w��F�o���#����ýmXýKv��fh}�:�>��&l����S֘�H���~��>��J����@��U��򘛾P   P   p����,��+�3������)��so𽲒�D%��ih}�Dd#�M�"�Gg���04�T8����-t�B��`S���E8�P   P   ��ɼS^<��c���xP��Y��d��FH �� ����Nv���jK�7������x#��>H{���1�����ی뽎���P   P   Cl�<�
�<�C;�������rĽ��GH �wo�qXý�������I�;8��<x�<~��<�]6<~�;8L*<���<P   P   z�=ySd=."=�G�9�%�
U���rĽg��-����ýAy��@���6�:D�=�Vg=bb�=�~�=��=�$�=��=P   P   �%�=݂�=��v=r��<���%�����Y������#������3����
=Z�w=��=O��=�:�=���=��=P   P   +��=�=�z�=|9v=p��<�F�9��輔xP�8���o���$P��2�\��9E��<�v=�a�=� �=~�=���=���=P   P   f��=2��=T{�=�z�=��v=,"=��C;�c���+���F���*�Gz���I;��=>v=d�=w��=�=�=;��=�C >P   P   1}>�?�=2��=�=݂�=ySd=�
�<X^<���,�� w�?wv�a+��l6�ŷ�<:d=��=�]�=���=���=�h>P   P   ���=���=:V�=���=���=I�J=mI~;P_�����,���@���+�q�[����;�J=��=��=0��=|v�=P   P   }v�=��=k��=�K�=���=�E�=��
<���J���ibѾz�о�>���HG�������<�\�=�7�=Y�=H��=P   P   1��=0�=�&�=�?�=���=?č=;�;�^������.��Mg�т�?�e��P�(�����$W�;΍=���=Y�=P   P   ��=���=>�=���=�:�=V.�=T��:���Z���9�ٿoH�?��j-ؿ</�������t;΍=�7�=P   P   ��=Lr�=�\�=4�=��=oR�=8{�;)���D�����!��o�^�����n�������U����=W�;�\�=P   P   �J=0Nj=3�g=��h=��l=��M=�C <k'���쾣���|7������:��-������mV6�������꾦����<P   P   G��;�ɺ<�Ĵ<I�<g �<���<YE�;<��,V������u ��_���x������Z��������=/�)������P   P   ��[�H�������Ἴ���'0��A��7�T�_�E�n
��/ؿ��n�&�������.����n�l-ؿ�P��HG�P   P   	q�
w�)p�52���g������Vmj�9o��l�˖��$�d�y��9��&���x���:��_���A��A�e��>��P   P   ��+�`�ƽ��½N�u������-��f���U(��ξ^���y���n��_�������o�qH��т�|�оP   P   ��@�z�`}����2/�rx8��`.�������G��<��ξ&�d��/ؿ�u ��|7��!�=�ٿRg�lbѾP   P   �,�=���@�Ϻ)��$N���c��:c�i�L�?�'�V���G�U(�͖��p
�������������1��Ŕ��P   P   ��𽹜ǽ,���x�)�I+Y�c?{������z���W�@�'����j���m�c�E�0V������D�`����J�P   P   P_�[x�@ý���o\N��r{�����ꉾ�z�k�L����-��Fo�E�T��<��v'�.������^�����P   P   [I~;�u��l�p����/��!d�Fڃ���������:c��`.����emj�^���D�;�C <�z�;�~�:��;��
<P   P   I�J=�`�<�X���{��(��89��!d��r{�g?{���c�wx8�������H0��r��<��M=kR�=R.�==č=�E�=P   P   ���=��k=�d�<Ŏ��hZ��(�� �/�r\N�M+Y��$N��2/�u��g�� ��J �<��l=��=�:�=���=���=P   P   ���=�B�={�h=駦<Ȏ���{���罶��|�)�Ժ)��+N�@2���Ἴ)�<��h={4�=���=�?�=�K�=P   P   :V�=���=�={�h=�d�<�X��r�p�
@ý3����@�j}����½?p�ҧ��dĴ<&�g=�\�=>�=�&�=j��=P   P   ���=k��=���=�B�=��k=�`�<�u��[x���ǽB��!z�i�ƽw�+H���ɺ<$Nj=Gr�=���=
0�=��=P   P   ���=>��=��=��=�;j=QD�<���0��O#��W�p�k�F�V��8"�!Ŀ�mA�ߊ�<kh=�y�=7�=.
�=P   P   /
�=)L�=���=)��=� �=�}<=��
��!���
M��g���ƾ�hƾ�\����J�uY��8�κ;=��=o��=��=P   P   7�=Ѷ�=���=���=c�={�l=|r��kN�@4��va
��G�؍`�z F�c	�PC��+��{ڹ��k=���=p��=P   P   �y�=R��=���=?��=Qt�=g�m=2��9�c���ʾ�IY�(ﵿ�쿎��5����W��,Ⱦ53���-:��k=��=P   P   kh=�5f=��a=�h=6}k=_�>=�a������ߗ�������F�.c�2LF�����E��a�߾53�xyڹ׺;=P   P   ���<S>�<\ă<\�<|�<��<����4�Ntɾ;��PW��ف�ԧ���� g��Q���E���,Ⱦ�*��7�P   P   [A��&ԼF�	�4�D���ʼoj��g�������W�b���������r������� g������W�PC��oY��P   P   Ŀ�:�DH����ѽo�н�ѷ�@��c��֦H�d������~9F�=������r������3LF�7���d	���J�P   P   �8"��~�����
1�):��0�x�t�����p��7�D���J�b�>�������ԧ�0c����| F��\��P   P   B�V���5��<P�`�u��߆�y����4t�z�M�K�2���R�E�þ�[^��꿀9F������ف���F���ۍ`��hƾP   P   n�k�*!Q��cv��A��I}���.���᪾���Bs��HM�s�f�F�þ9�D�����b�RW����,ﵿ�G��ƾP   P    �W��@Q�e��;�����ľǘ־�G־��þ� ��?g���HM���R��p��f���W�;��◊��IY�ya
��g��P   P   N#�BD6�(�v�������;�H�9:������̾� ���Bs�N�2���ۦH����Rtɾ⾞�ʾD4���
M�P   P   /������tP�+n��`ž;u꾁��������龆�þ��~�M�x��c��o����4Ὕ���c�rN彬!��P   P   ���0�����Iv��ޫ��׾�������;:���G־�᪾�4t�~�&@���j��$���g���9ds����
�P   P   SD�<��Ҽ�E���h1�}N���س��׾=u꾠H�˘־�.��}����0��ѷ��ʼ��<U�>=`�m=w�l=�}<=P   P   �;j=�J�<)��'Iҽ�;�~N���ޫ�cž��;��ľM}���߆�	):�}�нY���{�<,}k=Nt�=a�=� �=P   P   ��=�h=ݫ�<Q�(Iҽ�h1��Iv�-n������@����A��j�u�1���ѽK�;�<�h=<��=���=)��=P   P   ��=Cp�=
�b=۫�<,���E�����tP�.�v�i���cv��<P����SH��]�	�9ă<��a=���=���=���=P   P   >��=EO�=Cp�=�h=�J�<��Ҽ4�����ED6��@Q�1!Q���5��~�G�'Լ1>�<�5f=N��=϶�=(L�=P   P   J��=S�=\��=b�i=\��<�㮼�񤽞��.>_��`��Dg��,.����^�>��E%��>=��/��<�
g=b��=�Ƕ=P   P   �Ƕ=G�=��=t�=^b=5��<�"��H޽1�O���lⶾK����H��s�N��ܽQ�sȪ<�[_=!�=���=P   P   d��=�H�=Jz�=�l�=�^�=��'=���\�˽`>v��z׾�"�!')�y��;�վ��s���ɽ���ì%=��=!�=P   P   �
g=E�b=�c=J�i=��b=��(=Q�#��xҽ#j����	������o0���R~�J7�ٕ��Xн(Q0�Ǭ%=�[_=P   P   L��<q�<�?�<���<%~�<!{�<�a�dѽ�����mB�����X��N��������@�
7���Xн����Ȫ<P   P   =��,�����$�Y�꼨�����ǽ�B���A���п��0�3g�d�f�-P0��Ͽ�@�ٕ���ɽA�P   P   8%��9}���ݽQ��UJ۽�+�����9�ؽ\�r�RB�R��̕0�����ϖ����-P0�����K7���s��ܽP   P   6���&���C���W��W��B��#�v��a�K�8pԾ�}�'����f�sɖ��ϖ�e�f����R~�;�վn�N�P   P   ��^��o�m���(����!������o����k���Z����c(��E��=����f����5g��N�q0��z���H��P   P   (.�����Ї���ؾ/��eS��׾��Г�����j���R>'��E��(��Ε0���0��X�����#')�J���P   P   Ag��횧�ŚԾ���O��Z�Jl�{���PҾ���,���k���d(��}�R����п������"�lⶾP   P   �`������F߾V����*���9�)�9���)�8���ܾ����������;pԾUB��A��mB����z׾��P   P   +>_���u�Ծ'��w�2��rK��>T�z�J���1�8���PҾ�Г���Z�f�K�b�r��B������&j��c>v�2�O�P   P   ����<o�Q��������*�p�K�+^�T�]�{�J���)�}��򲵾�k�{��B�ؽ%�ǽmѽ yҽa�˽�H޽P   P   ���&��ߎ�j`پ�D�Ye:���T�,^��>T�,�9�Ll��׾�o��%�#��������a�ٮ#����"�P   P   }㮼��C����.�����Ze:�r�K��rK���9�Z�lS쾎���B�,����{�<��(=��'=5��<P   P   ^��<=Ｊ�ܽ�2X��Ӫ�/���D���*�z�2���*�R��7�쾪!���W�cJ۽���~�<��b=�^�=]b=P   P   c�i=�.�<x��H��2X����l`پ���*��Z������ؾ.�����W�a��:�e��<A�i=�l�=t�=P   P   [��=٩d=.H�<y����ܽ�C��ߎ�T���y�Ծ�F߾˚Ծׇ��s����C��ݽ��y?�<�c=Gz�=��=P   P   S�=1�=٩d=�.�<!=���&��<o���	���򚧾����o��&�I}��Y��Q�<;�b=�H�=F�=P   P   폔=��=�yX=j��<�x|�͓���.�e�ą��s����¾�鷾^y����e�������FY��R��<	YV="j�=P   P   #j�=HǊ=	=�K=p�<X-�YX������b��p���^��N>���&���b�����G����9�*��<�
H=R�|=P   P   YV=�2Z=)�W=�K=�h$=��<T�ļ�6ý��K��7��P|ܾ����۾�w��2�J���½�ȼt��<�� =�
H=P   P   i��<<�<��<�(�<���<$r8�C��p[T�nm̾1% ��nI�lI��q�90˾S�p7��p.E�~��<;��<P   P   !Y���ż��X/��g�u���"�����B����[�v�9PX������ı�*F���QW��+�|�Z�n7����ȼg�9�P   P   ���f,���н�5ϽJ����s���B������;xR����=>q�i ȿ����,�ǿ�~p��+�S���½�G��P   P   ���}�1���L���V�=�K�3�/����
�J_H��{ʾ>MW��ǿ`���x(�-��,�ǿ�QW�80˾-�J����P   P   �e�0=��zk��檲��A��2I�������a��F^�د��x��᛿+���h(��x(���+F���q��w���b�P   P   Xy��XZ���#��$�Y������?侀����헾i����Jپ��G���+��a�����ı�mI���۾�&��P   P   �鷾i��/����.���>�|�>�U�-�EK�0��Ӵ�+��x��§G�᛿��ǿk ȿ�����nI���J>��P   P   ��¾�a��^�)�`RT�c�s�W���r�9�R��(�k���Δ��+���Jپz��@MW�A>q�<PX�3% �P|ܾ�^��P   P   o���i��j~2�9�j�����~k��G(��C����h���0�l���Ӵ�k���گ���{ʾ���v�qm̾�7���p��P   P   ������澱�)�,�j�8���E ��*$�����������h��(�3�㾚헾�F^�O_H�@xR���[�s[T���K��b�P   P   )�e�^��g���T�)��M��ׄ��j>������C��<�R�GK�������a��
�����I���C���6ý���P   P   ��#���T澉/��dt��ۜ�I���؄��,$��I(����r�Y�-�@�������B������>r8�W�ļWX��P   P   }͓�pC1�$����m�z�?�I���ۜ�M��G ���k��]���>����8I��;�/��s����"����<��<X-�P   P   �x|������L����>w	�{�?��dt�)��;�������j�s��>�^���A��G�K�W�����u�x(�<�h$=p�<P   P   j��<����t�ϽE`W�����m��/��T�1�j�?�j�gRT���.��$����V��5Ͻ}/�����<�K=�K=P   P   �yX=���<��ݼt�Ͻ��L�&����T�j����)�o~2�d�)�5���#澁k����L��н!���<#�W=	=P   P   ��=�[=���<�������sC1�#��^�����$i���a��r��`Z��7=����1�v,����żտ�<�2Z=FǊ=P   P   �|E=�.=A��<l���u��b���_��K��D�Ҿ�9��|��{B����ҾƎ��oc`��I��Wy���!�!��<��,=P   P   ��,=v�-=��=�a�<P�ǻJD�l>ڽs�8�څ�qƪ�����v����Ǫ�R���?W9�zܽ=H���慢<�h=P   P   .��<���<��<�P�<�I7<����?��X׽2�;�d��w㮾6-��ʴ���7����;�͐ؽ��C�.�,�a@%<<P   P   }�!�ѢP�b�K�}�zv�����Ō��A����%�����žЖﾏ`ﾲž H��8�ᖽR���,���P   P   �Wy��T��^B��s͒�o�s�V A��k<���5A����Y���Q#���6�	#����ݍ�?��ᖽ��C��<H�P   P   }I��$!�b�1���0������"�ֽ��ӽ�z����E����)F��xz�\Zz�B�E�<����ݍ�8�ؽkܽP   P   bc`�G"��
l��'W���������I�\���5�í8�g���>�e�E��J�����<P��B�E���H����;�5W9�P   P   ����f�˾=��\����g�g�ɾ���������ALþ�M"���y�hy�����]Zz�	#��ž�7��L���P   P   �Ҿ�	��8*���B��K��B�_�(��r��TϾ^���?�������5���y��J���xz���6��`�Ǵ���Ǫ�P   P   qB����'�[�����R��v��_؃���X�aW%��:�.o���#����쾐M"�g�E��)F��Q#�Ж�3-��p���P   P   w���9�
]��啥�=�¿��Ϳ|)¿�J����}�2�6�>?��/o��@���CLþ�>�H���[�뾯�žu㮾����P   P   �9��1�9����U���)C�Ĵ��o�k��\ɸ�4���3�6��:�`������i��������&���d��mƪ�P   P   >�Ҿ�'��l�������T���,��w"�I������]ɸ���}�dW%��TϾ���ǭ8��z�7A���0�;�څ�P   P   �K��{	�B@[�'ҥ�f���[���.�ӄ.�J��n���J����X�s������5���ӽ$���A���X׽p�8�P   P   ��_�1�˾�U*�"ㄿ�ÿ�$�%�"���.��w"��o��)¿b؃�c�(�l�ɾP�\�+�ֽ�k<�Ό��?�h>ڽP   P   �b��Ԉ�s�zGC��ْ��ο�$��[��,�Ǵ���Ϳ{���B�g������d A�������FD�P   P   �u�]v ��\���Q���L��ْ���ÿj���T��0C�C�¿�R���K������������s��v���I7<N�ǻP   P   i�� ���H1�p����Q�|GC�#ㄿ*ҥ�����[���땥������B�a�/W����0�~͒����P�<�a�<P   P   @��<V�G������H1��\��u�U*�F@[��l�����]��%[��8*�H��l��l�1�jB����K���<��=P   P   �.=E��<W�G���^v ��Ԉ�5�˾~	��'�7�9���9��'��	�p�˾N"���$!��T���P����<r�-=P   P   $�<�&:<�[���?���ٽ�>C�Y���=�־�	��� ��)��� � 
�Ut׾�,���gD��@ܽ�C�q���5<P   P   �5<�8<#}�;��A��)�C���P�^Zn�+�,�Ⱦuf߾�w߾C+ɾpV���eo�`��aB����-�!cP���};P   P   R����������A��䨼w8%�*	��/2�y E��Y��q����媾s���ދ����E��_�tݜ���*�z'��cP�P   P   ߆C�C�S�ޡR���?��*(��B$�?�P�������8K�����t��r��DÈ�0�K�V���ᦽ�cW���*���-�P   P   �@ܽ�K��pJ�������ؽ���hP���̢�R
�25�`Æ��㮾�^��
ா	䆾�
6��齶ᦽkݜ�UB��P   P   �gD��Th�wJ}�ɚ|�"}f���A�;r��T ��Y��C4�nd������t龥
�p���∾�
6�R���_�W��P   P   �,��ڻ�twվ��޾�Ծ���Q����j���A��qH�ƻ��3���4��bU����p���䆾*�K���E��eo�P   P   Jt׾�
�m�$� �3��o3�y#�v���BԾ5S����������c��辯*�bU��
�	ாAÈ�؋��hV��P   P    
��:�˹j��ᇿ�����K����h���7�����tž���� ��㰽�辑4��u��^��r��n���9+ɾP   P   �� �We�/���V����ؿ�ؿ	���o����a�����U۾]���� ���c��3�������㮾t���媾�w߾P   P   �)�\��m���<��I/���#�&n������&����{��:&��U۾�������ǻ��od��`Æ�����l���mf߾P   P   �� �W���ſ4��B�Sje�1�d��NA����ÿ��{�����tž����qH��C4�25�8K��Y��%�ȾP   P   ��	�
e�����M(�W�T�Vߊ��&���)���R����&����a����8S����A��Y�T
����u E�&�P   P   7�־�9�hɚ�#��� C����%���ç��)���NA� ���r����7��BԾ��j��T ��̢����-2�XZn�P   P   V���F�	�[�j�tF�����Vf������%���&��7�d�+n�����h�z��V��Ar�nP��B�P�(	��
P�P   P   �>C�Aj���$�"��Piٿb�$��Vf� ��Yߊ�[je���#��ؿ�K��y#�����A�����B$�x8%�A���P   P   ��ٽvg��Tվq4��8��Qiٿ�� C�^�T�"�B�O/��ؿ�����o3��Ծ,}f���ؽ�*(��䨼�)�P   P   ��?�������|���޾q4�"��wF��)���R(�:��<��^����ᇿ�3���޾Ԛ|�������?���A���A�P   P   �[�i|Q������|��Tվ�$�_�j�kɚ�������ſ�m��6���ֹj�u�$�~wվ�J}�xJ��R����}�;P   P   �&:<��	�j|Q�����vg�Cj��H�	��9�e�
W�"\�ae��:��
�$ڻ��Th��K��S�S�����8<P   P   &�ټ�q�nyP����W��0~�/$����%U*���F�m<Q�@�F���*��q��쿾�}���	���R����P   P   ���"��Va���P�������އJ�0���¾_���@�?Q�<쾫�¾�撾1L��F�褽�bT�T��P   P   ��R�)�T�F,Q���P���f�%� �ؽB}�b\��E��Ҥ�����N��v���^�]�� �;	ܽa��Tl��bT�P   P   	��+Ž�pĽl,�����
q��H��SŽ�Y���4�5�a�~�o>~��pb���5�G��#�Ƚ�С�\���礽P   P   ��/�1�S9�V�0��*������ֽCĽ#�׽�	��A3��X�l�g��Y��04�M���۽�Ƚ1	ܽ�F�P   P   �}�����袾ʇ������s|�I�H�t��B��׵�/7&��vO���m�p�m��[P���'�J�B��� �&L�P   P   �쿾��#����f�����P\���S��Z�X��2��b1��N�Ms�������s��[P��04���5�S�]��撾P   P   �q��-���O�m(d���c�ruN�VR+�o��m%���Ɋ��]���U��l���������n�m��Y��pb�n�����¾P   P   ��*��~k����h���x弿�ڱ��P���h�D�'���쯡��py�E�d��l�Ms���m�g�g�f>~�G��
<�P   P   7�F�����8�ο���~���T�3̿�ِ��bC�{����E���py���U��N��vO�	�X�~�����9Q�P   P   d<Q��`������E�5�Kj�%��B�h���3��8��Pˢ���M�|�����]��b1�/7&��A3�/�a�Ҥ��@�P   P   ��F�Y��wn�9�Y��K�������W��	ڝ�
�V��n�Qˢ��bC����Ɋ��2�ص��	���4�E��V��P   P   U*��㒿����U�Y�*Ա��������������V��8���ِ�G�'�q%��_�X�D��#�׽�Y�b\��¾P   P   ��Gk���οW6�l���8����������ڝ���3�7̿�h�s���S��x��FĽSŽ?}� 0��P   P   +$��0�,�����,P���j�>���ϑ������W��K�h�X��P��[R+�U\��O�H���ֽI����ؽڇJ�P   P   ,~��o���O�,���C
�����@���8����������1�����ڱ�yuN�����s|����q��$����P   P   U��s���_���nd�����D
���j�q���1Ա�L��Xj��~��弿��c�l�����*�����f����P   P   �����0�ޚ��D���nd�.���.P�\6�^�Y�C�Y�N�5���q���w(d����ч��]�0�s,���P���P�P   P   nyP���ýV�8�ߚ��`����O�������ο����}n�	���C�ο�����O��#��袾[9��pĽM,Q�Xa�P   P   �q�oS���ý��0�t����o�3�,�Gk��㒿Y���`�������~k��-�$����8�1�4Ž1�T�$��P   P   �Ͻ��ӽzX轸���M���޾C��M�D��e�l�r�'f�&E��E���߾����v<O�wt��K齊"ԽP   P   �"Խ��ӽZ�нJ)ؽA��<m+��s�����&7ܾX���Q�Hh���gݾk���ռt��,�v� �y�ٽ�]ѽP   P   �K齾��ض�n3ؽ�&Ͻ>ླྀ6�V�9���t��b���ͮ��M�����=����uv��v;������9xѽv�ٽP   P   rt�A�j����h���ч߽#yֽR������3�q�U�̴j���j��V�YX5��k����=ڽ���r� �P   P   m<O��gi���r�2�h��{M�u�*�5Q
�8��Y"�5l���#��S$��V,�@�$�oi�<&��Z�罨�����,�P   P   ����ݞ���ľ��þm����"��gq�H�7�<�����������7��7�������7&���k��v;�ȼt�P   P   ��߾:/
�Om�N$�V��y	��ܾ���emq�:(1�Q�o��@	�Iu��<
���ji�PX5��uv�a���P   P   �E�K.J��u��[�����ps��H���	پ�ɕ�|�Q�ȯ!�FQ�l��Hu�7�:�$��V�4���[ݾP   P   E��኿���6Pۿ�9��5ڿQC����#B���;|��u�e��,)�FQ��@	�4���V,���j������P   P   �&f�򫯿_���cn*�I5H�_�G�� )��e��n����Fb�Y������v�e�ɯ!�n�����S$���j��M��@h�P   P   `�r��lǿN �6du��k��� ��
O���Xr����t!Ŀ�n�Z��=|��~�Q�Q�����#�h�U��ͮ��Q�P   P   �e�J^ǿ��-��?�����.2�+�����: ��l,+�u!Ŀ�Fb����ɕ�<(1����0l����3��b��S��P   P   F�D�P���sP ��M��:�H�2��6E�8�1�N� �< �����q���'B� 	پjmq�>��W"�����t�7ܾP   P   ?������%�����u����&�2�f�Z�fZ�:�1�	����Xr��e���������L�7�:��N��R�9�����P   P   �޾��I�bᶿ��*�
��$��Y�E�h�Z��6E�/��O��� )�WC���H��ܾnq�7Q
�#yֽ�6�{s�P   P   ���	���t�~}ۿ��H�_.��%��*�2�M�2�32�� ��i�G��5ڿps�~	��"��z�*�ԇ߽<�9m+�P   P   
�M��󳾳(��m�������H������?�����k��U5H��9鿚��\��s����{M�m����&Ͻ>��P   P   ���7ih���þ�W$��m���}ۿ��*�Ǟu��M���?��Fdu�mn*�BPۿ�[��N$���þ9�h���o3ؽI)ؽP   P   yX�&q��Ir���þ�(���t�fᶿ-���zP ���-�N �n�������u�Vm��ľ��r�n��ڶ�Z�нP   P   ��ӽ��&q�8ih��󳾥�	���I�����V���T^ǿ�lǿ�����኿U.J�A/
�垴��gi�E�����ӽP   P   �fv���n��Ma���b�JՃ�`S���T���@&��T���w��邿 7x���T���&�>v��6)���i���c��ea���n�P   P   ��n���n�^�\�h1F��|?�r�W��=�������ER��M��i�{��"��Y������R�X�B/@�[eF�J�\�P   P   �ea��l��sa�l?F�h*���Z*���O�	R����k������;��S���"����Q�Z,��+��+�ZeF�P   P   �c�Ty��,y��b��f?�����I
�!'
����8��2U���f��/g��7V�dK:�'���|���+�>/@�P   P   �i���Ж�g���P{��������V��)��	�6i����A9����4��0d����������T,�J�X�P   P   .)��~=о��Ȃ�/Ͼ����{G��
N���&m���rݽ�ڽ ޽��޽�ܽȤ���� ���Q����P   P   0v���f�Z.��K6�g�-��4�C}򾚤��k�����5�,n��tؽ�Ľ����i�ƽ�ܽ��ZK:�	"��N���P   P   ��&��\�w솿%����O���_Z��u$����T���JQ���� ۽�i��������޽)d��7V�J�����P   P   w�T�Y����˿�x��>B��/����ɿ>���2Q���7^��_b�-z�� ۽�Ľ��ݽ-���/g�1��r��P   P   7x�\���~A��F��fm�:�l�KND��d�����t�c��=��_b����tؽ�ڽ�����f�����i�P   P   �邿6|ܿxj7����������������א��4�x�ؿ����d��9^���JQ�,n�rݽ<9��2U�b����M�P   P   ��w�5gܿ�;H�kf��$���p/�>�.�0G�[���i�D�z�ؿ�t���T����5�&m������8���?R�P   P   �T��Y���_7�jp���o�)�Y�P�o���X����]����4�����2Q����n�����3i����R����P   P   �@&�����'��ϒ�Ÿ�C�Y�����VR����X�3G��א��d�B���u$�����N��	�'
���O����P   P   �T��q\���˿Z.F�Ga����/�/�p�����U�o�C�.�����SND���ɿ�_Z�J}�~G���)��I
�Z*��=��P   P   ]S��)��ӱ���~�� 	n�������/�G�Y�/�Y��p/�&���G�l��/��T���4�������V������n�W�P   P   HՃ��zϾ+�-��敿Z��"	n�Ka��ɸ�p�,�������fm�EB����n�-�/Ͼ�����f?�h*��|?�P   P   ��b��X���T�466��敿�~��_.F��ϒ�sp��vf�������F��x��-��K6�ς�S{���b�k?F�f1F�P   P   �Ma��x�gI���T�-�-�ձ����˿�'��_7�<H��j7��A���˿~솿Z.�(��k����,y��sa�\�\�P   P   ��n�^{l��x��X���zϾ+��u\�
����Y��@gܿB|ܿh���b���\��f��=о�Ж�Ty��l���n�P   P   m^��>���Ծ�Q��g����ľ�����(�buU���x�V)����x���U�r�)�� ��fž����-(�� �Ӿ���P   P   ���%��9-ھsر�gґ��=���Ę�@[��Җ�G��*7�7X�=	���II��4l��֘��s���>X��ޣپP   P   �Ӿ���oԾ�߱�Om���`��N���a�M��:��ɪ���~�����:桾���͑c��O��W`����>X��P   P   ,(��Roʾn�ʾi��Rԑ���_���1�HE�V&��<��U���d�Ae�n,V�$>�{!(�g� �t2��W`�q���P   P   ������Ǿ�Ҿ6�ǾN���������M�f���=�N� �����F�I!����S�<���[�c� ��O�Ҙ��P   P   �fžk0�9��>t��T�i$ľwm0`�R�$��+ ��ܽ�ѽP�Ͻ�н8�ӽh��9��t!(�c�-l��P   P   � �D( �x38��A�N�7�=�Fa�����(�����9�B��nϽ<V��l���`��3�ӽ�S�>����?I��P   P   h�)�m�a��Ŋ��К�y��	承N^_�@'�g��x����]Q������̽�6��l���н��b,V�0桾���P   P   w�U�;���Lп�����q��B��`Gο'��٬R���Om���R`�����̽:V��H�ϽA!�	Ae�|��5	�P   P   ��x�R�ÿ�BL��v���u�jmJ��1�Y����t����Թ��R`�����nϽ�ѽ�F���d��~��.X�P   P   O)��	=޿�:�(E��T����w��ŗ���Z��8�7���ڿ������Pm���]Q�B��ܽ����U�����#7�P   P   ��x�w#޿��K�b���G�Q6���5�F�����aPH���ڿ�t���z�����9��+ �J� �<�:��@��P   P   YuU��7ÿ��:��d���#���`��Ix�!�_�ą!�����;�7�\���ݬR�k��+���T�$��=�V&�M��ʖ�P   P   ��(�����%��wG�� l���`��ш�����#�_�I��Z���1�,��	@'����p0`�f��EE���a�;[��P   P   �����`��Ͽt9L�TQ���6�-�x��ш�Jx���5�͗��smJ�hGοV^_�Ma��z��M���1���N��Ę�P   P   �ľ����t���k���#w��w�� �6���`���`�Q6��w����u��B��承B�m$ľ������_��`��=��P   P   e���Jw�ͽ7�ê������#w�XQ��l��#��G�a���&�v��q�!y��U�7�U�O���Qԑ�Mm��dґ�P   P   �Q��O�ǾJM��@�Ī���k��z9L�}G��e��#b��3E��*BL������К��A�Bt�8�Ǿi���߱�pر�P   P   �Ծ{ʾVҾKM�Ͻ7��t���Ͽ*����:���K���:���Lп�Ŋ��38�=��"�Ҿn�ʾmԾ6-ھP   P   �>�����{ʾP�ǾMw������`������7ÿ�#޿=޿^�ÿD��y�a�K( �t0���ǾRoʾ���%��P   P   (�����t��D��L��� pݾ<� � �"��rI���h���t���h��I��#�N���ݾ02�����C��jt�P   P   �jt�e�t�=�P�����㾂H���e��	���>#�ڮ�Y��d�����	����)�������E��� ��P�P   P   ��C��T�5uD�4�����Cע�\���Qt�v燾�F��lR���e��ͫ��蝾O����_u�^��{��8�� �P   P   ����(�k)��P�����Ѣ�n=i���:���1��Y@��+U��dc��c��4V���A�g]3��e;���h�z��E��P   P   -2辗�
��~���
�ղ�-���:�t:�`�^`
����p�u�$(�P�9����e;�X������P   P   ��ݾ�1����$�����ݾD�����r�}�0���	�)�｠�佮�㽈�佻��o�6�`]3��_u�#���P   P   H�'�"��<�~E�s�;���!�l���~l���o����=�m�/5㽼˽�Ž ͽ���O���A�G������P   P   �#�@Y������=����*(W�G!��l������Q����-�R�ý�Ž���(�x4V�蝾x	�P   P   �I�|����ÿ���}���3�쿦8��5��JG�#��1_���*_��8��-ὺ˽���n��c�ë����P   P   ��h�(��M"���9�ԡ^���]��8����ڍ���Ze�]g����*_���.5㽚��~p��dc��e��\��P   P   ��t� �̿��(�/��<���Sz��[���n��Mf&�kɿq�]g�3_����Q�m�&�ｖ��+U�cR��Q��P   P   ��h�;n̿��6�7O���v ��!�� ��������4�kɿ [e�%�������=���	�[`
��Y@��F��Ԯ�P   P   �rI��ڴ�˪(��J�����02F��[�<YE�2�����Of&�ݍ��NG��l㾂o��~�0�`���1�q燾6#�P   P   �"�Ld�����M���r� ��VF���q�M�q�>YE����o�����9��K!��l����r�s:���:��Qt����P   P   9� ��rX�a�¿�x9�����"t!�J\���q��[��� �[���8��8��0(W�r���F����:�j=i�V���e��P   P   �oݾQ"��X�����^�d:��$t!��VF�62F��!�]z����]�>�����!��ݾ-���Ѣ�?ע�~H��P   P   
��4����;����a,���^�����v� �����v �H����^������y�;���Ӳ边�㾊����P   P   �L���
�����5E����!��x9�R����J��BO��8����9�����=��~E�&����
��P�1�����P   P   �D�v*)�ހ������;��X��f�¿���Ӫ(���6���(�V"��ÿ�����<�����~�h)�1uD�:�P�P   P   ��t�;�T�w*)���
�5��T"��rX�Qd���ڴ�En̿+�̿(������LY�.�"��1���
���(��T�b�t�P   P   X��%r�똵���q�c"�'���Ұ��-��o�3�q�L�m�V�� M��94�H��U���n��d�!�'%p�E�����P   P   ��[)�	�ƿ:$����1����ɼ����c�־�����*� ����׾Њ�����@�a0������iſP   P   H���+zǿ�\������:�S��0ܢ�5������������<��+e��j����2��"Ɇ�������Q08�����P   P   )%p��S�����j�q�&�1���tڜ�O�a�[4E�y�J��V\�|i�_�i��B]�}�K��F�F�a��������a0�P   P   e�!��F���U�RRG� s"�:��Ĵ��8�a��.�%��!�"�$+��B/�d�+�Ԧ#��; ��/�C�a����?�P   P   �n��Q����2��2�x������\��S��1D��=�
������j�����k��; ��F�Ɇ����P   P   �U����!�2�<�0�F��<<��R!�ľ��(ڻ��t��&�H��!�(����Z����	����Ϧ#�u�K��2��Ȋ��P   P   @�uF��_s�p����M��V5r���D�Sc�1�Ծ����CY���(����Zo�Y���j�^�+��B]�b����׾P   P   �94���}�B���7˿��ؿ�Vʿ�㦿`:{��1�Ƿ�[��H�e���,���������B/�U�i�"e�����P   P   � M�;!����#���K1�5�0�T���;߿U#��@/J�R�P��I�e���(�(���+�|i��<���*�P   P   b�V�w-��[x	�r�N����ؗ��R��J�L����Ҫ���S�S�\���CY��!�	���"��V\���� �P   P   h�L�e��_��w��&�����I������ҭt�X��Ҫ�B/J�ʷ���(�H��=�#��s�J��
�����P   P   h�3��ٚ�Z	�7{w�i���f���!��%�W��ԭt����X#��!�1�4�Ծ�t��2D��.�V4E����[�־P   P   (��L}�A3��N��4��s��I�2�`~2��%�����P�L��;߿f:{�Vc�+ڻ�S��5�a�J�a�2������P   P   ̰����E�Xͧ�r��*����:O"�K�2��!�P��R��Z���㦿��D�Ⱦ��\������pڜ�,ܢ��ɼ�P   P   "���K�!���r�#�ʿ�Z1�}��	��v��j���������=�0��Vʿ^5r��R!�����5����L���P   P   c"����n)<�?G��G�ؿ�Z1�!*��5��r����&������K1���ؿ�M���<<�x���r"�!�1��:���1�P   P   ��q��]G�ބ2��LF�@G��%�ʿu���N�B{w��w�~�N�,���7˿v���5�F��2�NRG�d�q����7$��P   P   阵����.V�ބ2�o)<���r�\ͧ�H3�Z	�_�cx	���%B���_s�7�<���2���U�����\���ƿP   P   #r�4$ȿ���]G����M�!��E�	L}��ٚ�n���-��D!����}�uF���!�S���F��S��(zǿX)�P   P   k�j���U�5��¿B|b��L�B�� �����q,���3���,�q�~;�<I������`�+��a��HU�P   P   JU�{xU�G_/��	��u������.ؾ���z�Ǿw�ݾ�A�t�'޾�'Ⱦ�����	׾`a�{Ӆ��{��4.�P   P   c���X/�[��Y�鿥�����*�ӧѾ�v��|p��@�����o��RT�������������թϾ�(������{�P   P   .���F����¿vw��1�*�a�Ҿ�E���Ch���f��zw����������Ex���g�_ah��o���о�(�|Ӆ�P   P   ��`�6뎿� �������b���T�Ѿ� ��hGY���H�<�P�h�]���c���^�%�Q�&�I���Y��o��ԩϾaa�P   P   ����=���X�,Y��>�+R���׾� ��Ig�vLH�-qE��*N�Q�U��ZV�@CO��G�$�I�[ah������	׾P   P   5I��G� ��o<�*G��n<�y� �S���� ���\����d�D�O�XyM��R��T�M�R�?CO�"�Q��g���������P   P   y;���.�{sT��k�Xak��S�U�-����ž%����t���[�ϬT��YT��T��ZV���^��Ex�����'ȾP   P   q���R��*��T��[��Sà��@����P�����ھS¡�����da�ЬT��R�P�U���c�����LT���'޾P   P   ��,�	�y�#�����/>��� ��߿`m����v��j*����Xצ�������[�YyM��*N�f�]�����o���t�P   P   ��3��O��;ο����a9��J�N�8�����*̿O����q1����T¡� �t�E�O�-qE�:�P��zw�����A�P   P   �q,�I9����ڿ�'(�+�n�s���eE�� >m�b�&�}�ؿP����j*���ھ'�����d�vLH���H���f�<���p�ݾP   P   ��zOy�fο�(���������6��%o���ǁ�c�&��*̿��v�����ž�\��Ig�fGY��Ch�yp��t�ǾP   P   ���AR����ڳ��n�!�����h��&o��>m����dm����P��� ��� ��� ���E���v������P   P   B���P.��͇��}�Y9�����'��������6��jE��S�8���߿�@��X�-�U�����׾O�Ѿ[�ҾͧѾ�.ؾP   P   �L��� �7�S�^���3��gJ�����!�����y���J��� �Xà��S�z� �)R���+�*���*����P   P   >|b���>�T<��8k�����3�Y9��n�Ĩ��6�n��a9�5>�b��_ak��n<�|�>�	�b�qw�������u��P   P   �¿я�_8Y��G��8k�`���}�޳��(��'(������T���k�*G�)Y����� �¿Q���	�P   P   3�������`8Y�T<�:�S��͇����nο��ڿ;ο,����*���sT��o<���X�� ����V��C_/�P   P   ��U��0����я���>��� ��P.��AR��Oy�O9���O���y���R�ƶ.�J� ���=�3뎿�F��X/�xxU�P   P   >���J)��:�k��t�߫���-�u:���r�sp�����>�Q��{�ﾨ��jV,��啿+����i�M���P   P   M������������/������L�����O'¾�D����;�ھ1?ھWXξ������������ J� ���(�-�@*��P   P   ��i�����3+k�¦/��Կ[f��������r)��ݣ�6G���v������)��H#���Բ��O�-�b��п)�-�P   P   .����/��P0�5:�����cf�lB�8���>ԑ��R��m�������Ѥ��f��ӧ��o���F��N�.�b����P   P   �啿�vſ�Cڿ��ƿ����0�L�4���q���鎾�������@�� ������Z#��s���@Ύ�F���O�� J�P   P   kV,�2�`�np���ab���-�~���T���=O��ƾ�����˶���ު�
���]�����r���n����Բ����P   P   ���5���<�Q�G�z�<�nL ������R��[��QK���ɔ�SO������}���]��Y#��ѧ��E#������P   P   s��m����4�^�G�y�G���4��K���頽��*��P���h��z��S`������
�������f���)������P   P   L��)��S���t�s倿�<t��Q�_�'�\J�L�˾���IĢ�s���{���ު�����Ѥ����PXξP   P   9�MNA�Q�	������n��<g��ju}��i?�&P�2׾��IĢ�i��TO��̶���@�������v��*?ھP   P   ��bLQ������)ÿ���E��]�)¿�Q��*O�gM�2׾���R����ɔ�������m��4G���ھP   P   ��S*Q��Й�{�ڿ�;�g�%�b�%�����mٿ����*O�'P�O�˾�*��RK��Ǿ������R��ݣ���;P   P   op���@�]���ڿ9��q@���P���?��g��mٿ�Q��j?�^J�렽�\��=O���鎾=ԑ�p)���D��P   P   �r��(���~���¿Z1��z@��b�I�b���?����,¿ou}�b�'��R��R����q��5�������K'¾P   P   p:������R��۝����6&��
Q��b���P�e�%�c�@g���Q��K�����x���0��hB��������P   P   �-��T ��4��lt�U���o��7&��z@��q@�k�%��E���n���<t���4�mL ���-�)�L��cf� [f���L�P   P   ۫��mb��<���G�1ǀ�V������\1�=��;���"���w倿}�G�y�<�ab�񟗿݉���Կ����P   P   �t�q7ǿ4���?�G���G��lt��۝���¿�ڿ��ڿ�)ÿ�� �t�c�G�P�G�꾂���ƿ/:���/��/�P   P   7�k�2�0�+lۿ5����<��4��R���~�]���Й�����Q��S���4��<�kp���Cڿ�P0�-+k�����P   P   I)��B��4�0�s7ǿmb��T �����(���@�Z*Q�jLQ�VNA�)�r��6��.�`��vſ��/���������P   P   j����c��	��C�7������VB�<����ܾ�A�\����w�� 6�������۾gX��$5@��X��ͦ5��v��_���P   P   `���4��?���,�^�%���Z3u��b�5�ξ�fľ}�ϾX�ھ,�ھ�8о�wľ�ξ��
�+Xq����+\�:���P   P   �v��_<���5���^����u͍����־���$�ľ��Ҿv'پ&Ӿ�žF޼�irԾZ���3��!>�+\�P   P   Ц5�a�]�Ks^�Ov7������͍�F�%�N߾(��[Ǿ�/ھ��羱�2�ھ��ǾQܿ��zݾ�#��3�����P   P   �X������D~�����ҹ��1u����I߾�h¾E�˾m�侦k��/+�\�����徚�̾�[¾�zݾ[��.Xq�P   P   '5@���}���o5��T���IB�b;�4pվ�s���{˾tQ�0�ؽ�J�������꾚�̾Pܿ�irԾ��
�P   P   gX��0���:�$�E���:����C����;U�����ž���������c�Hl���������ǾD޼��ξP   P   ��۾4��)���2'��3'�����@�K�ھ��¾Q�¾�+ؾp���',����c�J��]���2�ھ�ž�wľP   P   ����� �\!5�<8=���4�+g����⾋d;�5оNO�Q�(,���ٽ�0+���&Ӿ�8оP   P   �5��G��W57�,Y��Rn�.	n��CX�C6��)����׾y,־OO�r������0��k�����u'پ)�ھP   P   �w����LbL�P��i���i�����}~���J�d��I����׾�5о�+ؾ���wQ�p���/ھ��ҾV�ھP   P   X�������T������8��N���������������'$S�e����d;S�¾��ž�{˾G�˾[Ǿ%�ľ{�ϾP   P   �A侻]��0L�r���9b���}׿˟��*׿�Ӵ�������J��)��⾼�¾V����s���h¾(������fľP   P   �ܾћ���6�.	��$��q~׿Vg�H��*׿�����~�F6���L�ھ��;1pվ�I߾K߾�־3�ξP   P   8���{�����Q�X�K��T������Wg�Ο���������CX�.g��@��C��_;���A�%� ���b�P   P   �VB����{��[�4��n�-k��U���s~׿�}׿Q����i��3	n���4�������IB��1u��͍�p͍�S3u�P   P   ����O��ٻ:�H+'��=��n�K���$��=b���8���i���Rn�A8=��3'���:�J���ҹ�����������P   P   ?�7�,���~���<F�I+'�\�4�S�X�2	�u�������P�3Y�a!5��2'�!�E�i5�����Hv7��^�&�^�P   P   ��~b_�}a	�~���ۻ:�}�������6� 1L�ŤT�RbL�]57�	 �+���:���>~�Ds^��5��<���P   P   �c�����b_�/���Q�����|��ԛ��]�����L����6��/��{�}�����[�]�\<��2��P   P   ���a��#g��NG�zȿd�J�n���/�Ծ�Hؾ�"����V�1xؾ�ԾR���g>H�Sſ5�D��=������P   P   ����B��%���j�p�%�Q����M�az�ASܾ�뾉���7��n^��`ܾ^w����R��?��dn�pf��P   P   �=��������g�p��6�]A��b�0�>�����%V�a��p����������H���b.��E��Í�fn�P   P   9�D��o���o���F�����:���6;��	��������u"�|�.��.���"�4����$��n8��E��A��P   P   Sſ�u�	��z��'ȿ|��f�0����J��E>�rc4���J�xS��K��05���}��$��b.��R��P   P   k>H����nt��jF��c�J����7���:9�A��;��m[�fo�Lto�Md\�IP<�����H����P   P   T������u0�-;�a1�Vn�%�������_r3�w�Z�JTy������1z�Nd\��05�4����_w�P   P   �Ծ΂��~ ��
��
�Ջ �{��Ӿ=�پ������ ��I��n�'>������Nto��K���"�����`ܾP   P   /xؾf�޾_�����Q	��n�	���ܾ��վ%����
���,��=Q��n�LTy�ho�{S��.� �n^�P   P   �V��!�o@�����5���ZO�lK��q�@�⾌��Ql���,��I�z�Z��m[���J��.�q���7��P   P   ���M��� ��w'�o�:�	4B�9c:���&�����C���龍����
��� �br3�!;�vc4��u"�c�����P   P   �"�?-������4���Q�@d�d��TQ�=,3�����C��B��'�羚������D��H>����(V���P   P   �Hؾ8���W4�|�Z���x����	mx�Z�>,3�����q뾨�վ?�پę�;9�K�������CSܾP   P   /�Ծ�޾���M'���Q�D�x�W�����
mx��TQ���&�mK��ܾ�Ӿ�6�������	�>���az�P   P   l���s澺��O��ũ:��6d����W�����d�<c:�]O���{� ������a�0��6;�_�0��M�P   P   `�J����	� �
��� 1B��6d�F�x���x�@d�4B����n�ԋ �Rn�[�J�|���:��WA��M���P   P   �yȿ����{r1�8�
��	��Ʃ:���Q��Z���Q�s�:��5�S	�
�
�\1�dF���'ȿ����6�!�P   P    NG�1��(��@�;�8�
�
��P���M'�Z4��4��w'����«��
�-;��s���z���F�_�p�c�p�P   P   !g��f�p�!��(��|r1�
� ������������ �r@�c���~ ��u0�h���o����"���P   P   a��f���g�p�3��������u澁�޾:��C-���M���!�j�޾΂������{u��o����?��P   P   �����s��LR���	9��)��rC�-����e۾.%�΁��������V�4۾���S�@�� ����6��(��ϫ��P   P   Ы��#��¤��	�`�
^��P���M��������T�>����-Y���b3����s�|�D���M�]����P   P   �(�����M���h�`�U^
���Ԅ:������L�2��sG���O���G��q3��B�$��5H8�C������O�]�P   P   ��6�7^��^��8�����n����E��%�'�0���R���w��y������0�x���S��1�~�$�@_C�D���H���P   P   � ��]5��ZG�C��ƺ���l���+:���$��h8���f�EB��] ������������h�{}9��$�7H8�w�|�P   P   W�@�#{s��7�����G�u�R�B�g���J�i�/��f�����C����οQ3Ͽ"8���ܗ��h��1�&�����P   P   ������N��T�%�@���oa��?i �vW�	Q��Z��އ��B�ڿ�
�e�ۿ#8������S��B�d3�P   P   6۾O\Ͼ�g׾G����]Y׾��ξ��ؾ����l0���t��y��3�Ϳk��
�S3Ͽ ���4�x��q3���P   P   �V�V�ž�ÿ�x�þw�ƾdxþ]����Cþ��߾��0-D�4������4�ͿD�ڿ��ο����������G�/Y�P   P   ���hѾoȾ�̾9Ҿ�Ѿ��˾K]ƾWξ*����.�K�5����y��ᇸ�F��a ���y����O���P   P   �����Dܾ��־�v�L�쾡�Z�n�޾]YԾz�ؾW������2-D�ít��Z������IB���w��sG�A��P   P   ҁ�e.ܾ !ݾ*�	3��k	��C	�-����߀ھ{�ؾ+����l0�Q��f���f���R�Q�2�X�P   P   2%㾩=ѾT�־�l��4Y�����2�	��^YԾXξ��߾���xW�m�/��h8�+�0�������P   P   �e۾��žZFȾ�Q��'�dZ�ϣ����.��p�޾M]ƾ�Cþ��ؾ?i ��J���$��%������P   P   -����оQ翾��̾~���p	��+�ϣ����C	�]� �˾^�����ξka��c���+:���E�҄:�L��P   P   oC���]Cؾ�ľ[EҾ�8��p	�eZ�5Y��k	����Ѿexþ[Y׾��K�B��l���n����M���P   P   �)��gv����iH⾣Ǿ[EҾ���'����3�O��	9Ҿx�ƾ��@�<�u��������O^
�^��P   P   �	9�UL���|���&�jH��ľ��̾�Qྌl�,v��̾y�þD��O�%�����7���8�a�`��`�P   P   KR��/"`��h��|�����^CؾQ翾ZFȾU�־!ݾ��־oȾ�ÿ��g׾I���7��TG��^�I�������P   P   �s��֬��1"`�XL��gv����о��ž�=Ѿe.ܾ�Dܾ�hѾV�žM\Ͼ���{s�T5��7^����#��P   P   賩�ԛ�Oqn��h�be����.�Co��d�@u���i�����@���O���3�,�D��OT��Vl� /��P   P   /����������N3�6�ɿ�)d�JM ��p��i&� >���M���M�]x>���&��k��'���`��>ƿ"�0�$���P   P   �Vl�1����m��3�AD޿��$�<���2��N���y�
!���m���}����z���O�D�2��4;��	���Oڿ$�0�P   P   ST�mW0���0�����{ɿ������G���D��Do��ș��i���pԿ��Կ�^��]䚿��p��WE�,7F��	���>ƿP   P   H���w��n�Կ[�¿�똿.�c�W<��gD�M7{���� ��l
����
���q����}��WE��4;���`�P   P   7�,��UL�uf�2#g��M�b'.�TN�mv1�^�m� u��o���p78��8�$i �w���r�����p�F�2��'�P   P   ��h~������>x�F�����u��WL����ĸ⿟j���F��#X�46H�%i ���_䚿��O��k�P   P   �O�Q¾�봾���g�����������#��eu�ސ��-r�<�6��EW�$X��8��
��^����z���&�P   P   C������ϟ��7��Z�������V���R������v:�II��ӗп,��>�6���F�u78�
����Կ�}��bx>�P   P   ���Tξr量����*玾�~���+��WB��4�ɾ�T
��I�&��ԗп/r��j���q
��pԿ�m����M�P   P   m���2ھ�y���̟�f���H��O����松K:��V9վ*"��I�KI��ᐺ�ɸ�w��(���i��!���M�P   P   ��Rھ����D�������9䧾ǆ���s���y��N)��W9վ�T
�x:��eu����&u������ș��y�'>�P   P   Du�y(ξ�g��L���`���K~�����갾c@���y��L:��5�ɾ������#�WL�d�m�U7{��Do� �N��i&�P   P   $d�`����᥾�ɟ�ѣ��Џ��n��Q۸�갾�s���松XB���R�����v��ov1��gD���D���2��p�P   P   Fo����¾���㫔��������ON��n�����Ȇ��P����+��V��������SN�U<���G�$�<�JM �P   P   ��.����2ܵ�4���<=��ݸ�����я��L~��;䧾�H���~������g��@���\'.�'�c��������)d�P   P   _e��1�N��:�I��s4��<=������ң��a�������f��+玾Y����:x���M��똿�{ɿ9D޿0�ɿP   P   �h��ÿb�h�>�	�I��4���⫔��ɟ�L���D����̟������7����� ��(#g�R�¿����3��N3�P   P   Lqn�2��ֿc�h��:�1ܵ�����᥾�g�������y��q量ϟ��봾��uf�e�Կ��0���m����P   P   ԛ�t���2��ÿ3�N������¾\���t(ξNھ�2ھTξ�����P¾b~���UL��w��hW0�/������P   P   8�n��Y��%"���ƿ��e�O����� M����!�*��32�A+�FQ���������-�C�b��ÿۅ ���X�P   P   ��X��+Y�xA3��i�v���A@�E� �k�,���O�Sv�<_��������v���P�N-��7 ��F>�������1�P   P   ݅ ���1���!�q�k��,[��<���Q����s|��%ʿ2�ֿB�ʿ"���������R�C�;���X�H������P   P   
�ÿC��"��ſ�ԑ���Z��dF�](h��ߝ�1ۿ����#�V)$�l��)\ݿ[��� �i��IF���X���P   P   H�b����Ȓ�;숿�d��?�	D;�+jg��-����=3��Af��|���g��M5�/����c��!�i�E�;��F>�P   P   �-��=�z�+���+�K���z��?���O�]�������bB�Vr��oѩ��������:�E�1���]�����R��7 �P   P   ����ThؾBbҾ��Ӿ�pҾѷ׾�2��Pj*�P����DؿlV1�꜊�&P��$���
������M5�-\ݿ����Q-�P   P   ���p5���E��gS��������b��7��׬K�����W�+mb�2���}��&���������g�o��&�����P�P   P   JQ���Ǿ}|���=k��C\�E0i�S���#þ�?��p��0ſz��c3w�4��*P��tѩ��|�\)$�I�ʿ��v�P   P   A+�S�ݾ�ۘ��j��[M�DCL�<$g�FR��P|׾y]&�õ��Iѿ{��/mb��[r���Af���#�:�ֿ����P   P   �32�q��+��	�{�}�V�EK�z_T��w��頾� 澈!-�õ���0ſ�W�rV1��bB��=3����/ʿB_��P   P   (�*��쾊b��zƄ��2d�\NU�y_T��;a�� ���륾� �z]&��p�����Dؿ���9���1ۿ||��^v�P   P   ���]Iݾ#���Ǆ�j���]��3Z�B)\��f�� ���頾R|׾�?�ڬK�T���b���$��ߝ������O�P   P   M�a�Ǿ�՘��|�/wd���]�[o]���\�B)\��;a��w�GR���#þ9��Sj*���O�2jg�e(h���Q�q�,�P   P   ���ꓽ������Ik�R)W��V�>�Z�[o]��3Z�z_T�|_T�>$g�T���b���2���?�
D;��dF��<�H� �P   P   P����پd���_l�وN��L��V���]���]�\NU�EK�DCL�D0i����ͷ׾�z��?���Z�,[��A@�P   P   ��e�1� �AԾ�g���/^�׈N�Q)W�-wd�j��2d�}�V��[M��C\� ���pҾF���d�~ԑ�f��s��P   P   ��ƿ庉�3-��Qվ�g���_l��Ik��|��Ǆ�xƄ��{��j��=k�dS����Ӿ|�+�6숿��ſi�i�P   P   �%"����R��3-�AԾb�������՘����b��+���ۘ�{|���E��;bҾt�+��Ȓ��"���!�tA3�P   P   �Y���2����溉�2� ���پ哽�Z�ǾUIݾ��k��M�ݾ��Ǿl5��Ohؾ�=���C쿟�1��+Y�P   P   R>	������&����v���$��| � ���N�2�H�K��uU��L�Ɓ3�ќ�?��Բ��hN#��t��T��E_��P   P   G_���!��tͿ����J��< � �!���D�o;{�Nq��n~������)��J�|���E�u�!�1c���H�l`��^;˿P   P   �T��rʿ����呿X�Y�T�3��;�/�p��ӥ��(޿v�G���
���߿N^��;�r��~<��3��pW�m`��P   P   �t�'��6r���u��*J���3��tE�ݲ��~�ǿ��gJ�usr�<s��6L�����Qʿ"K��S�F��3���H�P   P   kN#�uu3�w/<��/4�$��P���:�M0��_Կ�,��!���������x���4��r
0�]ؿ#K��<�3c�P   P   ٲ�� �����_�(���y�����n�]�ſ��+�"e�������{0��=������s
0��Qʿ>�r�w�!�P   P   ?�� ����٣��ڝ�F��H���,����kA�����o�TL���~������-�2<� >���4�����Q^����E�P   P   ՜�����d����c��b�ϱ����������u�rٿ��E�/E��>��E�,��-�~0�x��7L���߿Q�|�P   P   ́3��h׾@����9G�|"0��wD�PV��?LѾ�.�7��u��d?k����@�������'���&<s��
�.��P   P   �L�&��Y瘾"NM��n!�� �0�H�j��NI�
�E�u&��o��f?k�3E���~����������sr�N������P   P   �uU�S��̧�+_���%����#��X�w{���� ���N�v&��v����E�YL��*e���!��gJ� v�w~��P   P   Q�K�T��3����%l���.�<��s���+��Ce��+���� ��E�7��wٿ�o���+�"�,�&���(޿Vq��P   P   W�2�)��� ����0l���2����Tq�{��	�.��Ce�x{��PI.��u�����e�ſ_Կ��ǿ�ӥ�|;{�P   P   �D
׾P٘��]_��9/����:���,�{���+��X��j��ALѾ����kA��n�R0��㲅�:�p���D�P   P   " ��Ѷ��������M�Ѯ&�������9��Tq�t��#�1�H�QV������/���	����:��tE��;�&�!�P   P   �| ��`���1����H��"�������������;������ ��wD�ϱ��G����y���P���3�T�3��< �P   P   ��$�`	�K����e�G}2��"�Ϯ&��9/���2���.���%��n!�z"0��b�F��#��$��*J�U�Y��J�P   P   ��v�]5�X�e����e���H���M��]_��0l��%l�&_�NM��9G��c��ڝ�W��/4��u��呿���P   P   �&���[����=�X�K���1������J٘�����-���̧�U瘾<���`����٣����q/<�1r�����pͿP   P   ������˿�[��]5�_	�`��ʶ��;
׾���N��O�����h׾����������pu3�$��nʿ�!��P   P   �Y��E�{�{�I�6��B_�RK߾[� �d|"�^,I��Yh�ڐt���h�YJ�DO#�{b��1߾f��x?��H�|�z�P   P   ~�z��4{���Y���,�����+"�,�W��Տ�]&����˿�#̿���䐿I�Y��!#�/��2�z+��aX�P   P   �H��lU�n�H�J�,�������CR;���+��B��d�'���5�Ac(�}$��Zÿo$����<�p����z+�P   P   z?��| ��� �������L��ZD�������47��@������G=������9�_������l�F�q���2�P   P   k��z~�Z�����a������:���������Z��-���(��b��b���^���p_��< �������<�1�P   P   �1߾��������&g��H��=ܾu �~��ʚ��Y�������pRC�2D��d �M����p_�b��q$���!#�P   P   ~b�J���o��6	k�����즾������S�-���U�3��u�������W��nn���Y��d ��^���9��ZÿN�Y�P   P   HO#��=��7kv�P<�O�:�f�q��4��+��T��`������������@�;4m��nn�2D��b��#����$��䐿P   P   `J��T羸���%�3�ue�CQ0����
�߾fC������#"��'��q�	���@���W�wRC�b�O=��Ic(�	��P   P   ��h��"��Q���dB����[
�8�<�S���w�z�`�t�ĿBA/��'������������(��Ꝣ���5��#̿P   P   �t����4��gRW��1�����h9P�/�������)l�u�Ŀ�#"������u�������-���@��o�'���˿P   P   �Yh�����	���ke����O齌�����`]��{�����|�`�����d��\�3��Y��Z�@7�J��g&��P   P   i,I����D��O}e��n��%齼�Ͻ��佺���`]�0����w�
fC�T��4���Ԛ��������+���Տ�P   P   l|"�ǳ�#/����W�wS�f��-�ʽv�Ƚ�����j9P�U���߾/����S�������ů������7�W�P   P   a� �nۿ�L��C�m;�]�뽱vҽ,�ʽ��Ͻ����:�<�����4������y ��:��ZD�KR;��+"�P   P   YK߾p詾Gw� 5�B��ߗ��[��b���%�O齏���[
�CQ0�h�q��즾?ܾ���L������P   P   E_�8�����!>�D	�@��i;�sS��n�����1���se�M�:����G��_�꾪������P   P   6����辫!����m��!>�5�
C���W�G}e��ke�`RW��dB�!�3�M<�1	k�"g��������G�,���,�P   P   z�I��!�۾꾪!����Gw�F��/��<���	���4���Q������0kv�l��󖤾T�辋� �j�H���Y�P   P   C�{��V��!����5��j詾eۿ���澭��������"��T��=��F�������u~澞| ��lU��4{�P   P   v��L����پ�|���l��otƾf3 �-�)��V��y�o����<z��0W��*�y� ��/Ǿ�2��hx��:�ؾ�b��P   P   �b������6���Ͼ�ʾ 4� �*a��䙿�ÿ;�޿rV߿�Ŀ2���_c�~z!����;�ʾξG��P   P   <�ؾ'P߾�پ��ξ�վ�����7�?=����Ͽ ����:�{�L�[<��S�g9ҿ����:��j}վξP   P   kx���]���v���p����ɾ���b:@�U���-���:K���l����i��付�Y�N�� �ў��>9C��=�ʾP   P    3���7����Oȓ� ì��뾏z6�
4��Q:��pt����8���Q#�cG�����
�z��t
�Ҟ���:����P   P   �/ǾZ)��JIc��cb�?����þ��������`��5�r����[45�'`�Fa���7�����z�� �����z!�P   P   |� �k���X@Q��I3�vcN�~2��j��&�\��˿�WG�L�����3�i�v��z���?y���7�����^�N�l9ҿ�_c�P   P   �*��p���d�(� �N�m_�봺��5%�q���������
��9I]������z��Ka�hG�뻘��S�"2��P   P   �0W����pψ��S(��3��{$�}d��E��X�O�@v���u4������;I]�n�v�.`��Q#��i��e<�%�ĿP   P   �<z����Ģ��>��d�'� �ַ8�f蜾k�	�+q��ֿ�nD��������3�b45�@��x�����L�}V߿P   P   v���m����zkW����&�޽s8���O�F6���a�&�}��ֿ�u4�����U��������������:�H�޿P   P   �y�\������
g��2��Խ$ѽHw�A^��w���a�+q�Dv����XG�C�r��pt��:K�*���ÿP   P   �V��c�'趾5"g�[��=ӽ9��jMν��A^�G6��l�	�\�O�u���
�˿�`��Y:�<��
�Ͽ�䙿P   P   7�)�}��X�����W�����&Խ>����֮�jMνHw��O�i蜾I���5%�.�\�����4��]���G=��*a�P   P   m3 �?�������~i?���	���ֽ4ι�<���8��#ѽs8�ط8��d��ﴺ�q������z6�j:@���7�� �P   P   xtƾ@_��[2e�8�)��R������ֽ�&Խ�=ӽ�Խ$�޽'� ��{$�q_��2�� �þ�뾭�����)4�P   P   �l������Z�R�o�"���	��R���	����V��2�����d��3�N�wcN�@���ì���ɾ�վ�ʾP   P   �|���3���Ke���5�l�"�2�)�ui?���W�,"g�g�rkW���>��S(�%� ��I3��cb�Nȓ��p����ξ�ϾP   P   ��پ����
���Ke�T�R�Q2e�����O���趾�������Ģ�lψ�޾d�T@Q�FIc����v���پ5��P   P   �L��vྀ����3������9_��5���p�ﾜc�T��f��������p��g���W)���7���]��$P߾����P   P   �{~���v��*h�hh�V���@��`r��Ё'�h�U�#z��1����z���V�P�(��S���|�����>�g��dg��9v�P   P   �9v�%vv�Ys�C|~������;Ѿ���=]�K�����¿��޿!߿{ Ŀc��F�_��r�BӾKn���~���r�P   P   �dg��b��Gg���}��"��k�㾣}.�����y̿���69���J��c:���9;Ͽ�
����0��}�酠��~�P   P   @�g�+2K���J�l]f�b���y��= 6��͕�����#�F����uǸ�왹�:���qJ��\��Z���Al9��}�Ln��P   P   �����C��-�#B��v��U$Ͼ�1-��'��T��m�F ����� �#B�����-�s��F�[�����0�BӾP   P   �|��a�[�--!�7����W��R������b������l�@����]0�w[���\��3�e���/�s��\���
���r�P   P   �S��S�����-��D�^M*��ꈾW�]�X�^�ȿ-(C������'/��,q�������s��3������qJ�>;ϿK�_�P   P   U�(�Z���C�S�T��
�,�M����2#��Ҕ�A��ˏ�<���X�����������\�(B�@����h��P   P   ��V�9��a����o���@��3ǀ�F��AVO��ȼ��2�5D���F��X��,q�w[�� ������c:�� ĿP   P   ��z���(!���;�aX�������C5����H�	���q�6�ֿ��B�7D��?���'/��]0�'���Ǹ���J�!߿P   P   �1������߷�
X�L	�";߽�]�`�O�Lϰ�+�0�~�8�ֿ�2��ˏ�����M���T �� ���69���޿P   P   0z�n���쿾��i��t��5ܽ;)ٽ���at`�R���,���q��ȼ�#A�6(C��l��m�2�F�	���¿P   P   t�U��������W�i�GN�w)�B�Ž۽���bt`�Nϰ�J�	�EVO��Ҕ�e�ȿ���\�
����y̿T���P   P   ځ'��ҡ��9X�v���ὡ½�7��۽���b�O����K��2#�e�X�c���'���͕����=]�P   P   nr��ē��� ��<��
��޽(�Ƚ�½A�Ž;)ٽ�]��C5�5ǀ����_񾮋��1-�F 6��}.����P   P   �@����K�S���O ��C� �޽��s)��5ܽ ;߽����B��1�M��ꈾ�R��]$Ͼ���v���;ѾP   P   \����[��p.��mK��M ��
�q��AN��t�I	�\X��n����
�aM*���W��v��g����"������P   P   nh�IxD���"��a����<��9X�L�i���i�
X��;���
T��D�8��#B�o]f���}�I|~�P   P   �*h��ZL��/��"��p.�@�S�� ���ҡ���쿾�߷�"!���a��>�S���-�+-!�~�-���J��Gg�Ys�P   P   ��v��d��ZL�DxD���[���������ٟ�f�������1�U���P���]�[���C�)2K��b�%vv�P   P   �yٽ�tݽ������R�1�����w���GG�0i�|jv���i�}H������ᣜ���S��{�?��a;ݽP   P   a;ݽvݽ����͆!�t7l��������K�+L�������ʿ�)˿�!�������N����H���n�[�"�w���P   P   @��"ٽJ�.� ��du�i8ž�5�U�v�Ŷ���x�E'#���1��*$�^��V=���Mz��� �XWȾ��x�[�"�P   P   �{�?ཷ߽i��j�3�ľ�$�Q�����ܿ��,��z�Q������<}���/�'�O����(�YWȾ�n�P   P   ��S����o�ս���<O��
��P�yh��>}�
XJ��E������t}�BQ��o���CCO�~"�P����� ��H��P   P   䣜��C0�ɩ潵�H,��m��:	���s��ڿoI�����J��j�6���7�5� ���ECO�'��Mz���P   P   ��*y��R۽{��z{q��ܾ��G�uN��x�)��ͥ�}��{�H�J=_�P�J�5�r�����/�Z=���N�P   P   ���mL���#>��C򽆤)8��y�����|و��j���^s������^4�J�]�M=_���7�JQ���<}�b������P   P   %}H��u�kz���ʡ�l���%q��\ؾ�hA�"���&������]���^4��H�o�6�z}�$���+$��!��P   P   ��i�< �
!���97����:Y��11�zN����	sa���ÿ�,+������������Q������Z����1��)˿P   P   �jv�ϑ�2����	Y�z��$w��IM��=Q��ª�����m���ÿ)���^s��ͥ������E���z�O'#���ʿP   P   !0i�^d�]ӹ���m�7�%��K�!���!���d��̲���sa�&���k���)�zI�XJ���,��x����P   P   �GG����I��[�m��-����"����iT(���d��ª����hA��و�|N��)�ڿL}���ܿж��3L��P   P   ����c߾����bY�T&��6�@��N�
����!��=Q�}N���\ؾ�����G���s��h��Y���c�v��K�P   P   �ᾭD��r\y��|7�����d�*�	�@��"��"��JM�41��%q��y���ܾ@	�X��$��5���P   P   1��t�w�C�=� ��� ������d��6�����K�#w��<Y��n���)8��{q��m���
��=�ľt8ž����P   P   �R�r�/����2���Q�� ����O&��-�3�%�w�����ɡ潊����O,�FO��j�eu��7l�P   P   ������w轼߽+�����|7�XY�Q�m�|�m��	Y��97����C�R۽�佪��i�5� �Ն!�P   P   ��F$��׽�w轝��9�=�d\y�����I��Tӹ�+���!��cz��#>��ǩ�q�ս�߽J����P   P   �tݽ�ڽA$���h�/�d�w��D���c߾��Wd�ȑ�6 ��u�gL��#y��C0����?�$ٽxݽP   P   Z���:��,7_��载�!������¾ek�f]-��`J�ԔU��	K�"s.�m���ľ���f�"��ο���`��N�P   P   �N�h�o�`���ʽ��4�)�Q���i/�u8o�Kŕ� ��|o�������oq�u1�	��-��v�7�?νd�P   P   ��`��>&�	N]���ɽ��;�^���h��8R�������ҿ���I=�	����Կ����JiU�b�	�蝧���?�?νP   P   �ο�z�_�]��_���Y3�z ��z
��vf��3������:���`���a�A�<�X�	�+w��9�j�"��靧�w�7�P   P   h�"�97�� �s�B5���_�7��1y�I�e�t+���9��gp�cϤ�C��y~����t�,���ÿ:�j�c�	��-��P   P   ������K���Ě���a~�{L���O�����b�u��� ��x����4�������o��-��-w��MiU��P   P   ��ľ�4Q�SD��ꣽf�ڽ}/J�`B���,�tV��ę�B<m�����u
�Uc���������t�[�	�����u1�P   P   q���E��1�#�7�˽NoȽ:���������i��Ϳ1[6�ac���u���w�Vc��4��~~��G�<���Կ�oq�P   P   (s.���ƾ�b�;�	�TܽB��Y�����j_(�����Q��5�Y������u���u
�����J����a�������P   P   �	K�V�P��e38�OA�ׂ	�d�2�z��]7辜�C�;�����8�Y�ec������� ��lϤ���`�P=��o��P   P   ޔU�����ϧ�B�d�%4�l&���0��]������ ��;N�<���"Q��6[6�L<m�|���gp�$�:����	��P   P   �`J�����z���;��ѧX�V�M�z�L��wT���x�q<��� ���C�����%�Ϳə�&b��9������ҿSŕ�P   P   p]-�82�+|��B#���Wg���j��o���h���b���x�����`7�n_(��i�zV������~+���3�������8o�P   P   mk�6�žϏ��ad�ِX�5�j�	���~���h��wT��]�}���������,���O�T�e��vf��8R�j/�P   P   ��¾:���(a��8�WR4�q[N��Dp�
���o�{�L���0�g�2�"�Y�����gB���L�8y��
�p�`��P   P   ���ߢO�+#�[6
��%��U'�p[N�4�j���j�V�M�l&�ق	�E�?��/J��a~�7��� ��h���3�P   P   �!�V������ͽ��߽�%�SR4�ՐX�|Wg�ϧX�%4�OA�UܽSoȽo�ڽ"��_��Y3��;���4�P   P   �载���� ���@	����ͽV6
��8�ad�>#���;��<�d�a38�8�	�5�˽�ꣽ�Ě�L5��
`����ɽ��ʽP   P   ;7_�TI`��kw�������+#��(a�Ϗ�#|���z���ϧ�~P���b�-�#�ODὠK��'�s�]�N]��`�P   P   ?���#'�KI`������U�ѢO�:��*�ž,2𾍳����M���ƾ�E���4Q���87��}�_��>&�h�P   P   �o<s�<�MJ���O�Vp�sI�U`��p�۾�
�k$��_-���$�=����ݾ���}�K����V�S��'R�q�<P   P   z�<��<��=��_��*��m�@V��[���>��j��!���e��� l���?�m[�'¾� q�]���,f��J�P   P   �'R��ǟ:��C��>^�����怾u�ؾ�e'��o�|����Ӿ�̿Pӿ�2��n�r���)���ܾ��� 
��,f�P   P   W�S�)<~���s�cLK�6����Y�����˦6�����ſ�n��?����]��oȿwˌ�:���� ���_��P   P   ��潝E;��ļ%�3�.�޽*j��J׾�5��,��3�ݿ����^J�U^��L�7 ����.3��:���ܾ� q�P   P   ��K�𾽌45�*�0�������D��c��!�%��]���ܿE�(��qn�)^��o#���q�6,����yˌ���)�+¾P   P   ����L#�,X���^������+��ʘ��
���k��ÿw<�"�l��ܞ��c��ߩ���q� 7 �!oȿs�r�p[�P   P   ��ݾ��v�S~������觽w���m��\־�9��<������V�F�.����T���c��q#���L�`��6����?�P   P   B���ç�\�J��2	��
�#��`�C�G����	��vd�6�0���RY�/����ܞ�-^��U^����Vӿ�� l�P   P   ��$��$ξT3����M�g�5�[4���H����B�ƾ�\��~~�2ƿ1��Y�F�)�l��qn��^J��?�̿�e��P   P   �_-�����+��5e�������������Y�����^�ܾR�'��~~�9򹿍���|<�L�(�����n��Ӿ��!��P   P   k$��C�"E��᎟�&��ɮ��/'���Q���W�����_�ܾ�\��vd��<���ÿ(�ܿ>�ݿ�ſ�����j�P   P   �
�J;�����N���μ��l�����&��=4���W�����F�ƾ�	��9���k��]���,�������o��>�P   P   }�۾걦�L|���Ј������%�����'���Q���Y��	���K����\־�
�)�%��5�Ԧ6��e'�c��P   P   ``��x�t�yI�ȱL�4����(�����������1'��������H�f�C�
�m��ʘ��c���J׾��ᾂ�ؾLV��P   P   �I�:�!�*������5����(���%��l�ˮ������[4�'��}���+���D�9j��Y���怾�m�P   P   kp�-A���5���竽����5�3��������μ�'�����i�5��
��觽��������@�޽L������*�P   P   ��O���9�x�6���b�{竽���±L��Ј��N��ߎ��4e����M��2	������^�7�0�8�3�|LK��>^� �_�P   P   �MJ��a~��mʼm�6��5��!��nI�G|������E���+��Q3��W�J�P~�)X���45���ļžs���C��=�P   P   ^�<�:�a~���9�A��.�!�h�t�ᱦ��I;{C価�侾$ξ�ç���v��L#��ﾽ�E;�:<~��Ɵ:��<P   P   6Y9=Q2!=�<9 W�é���g�,g� ���fؾ�4���������پ\���-j���������d��]�<{ =P   P   { =�^!=��<_x��N��~v&��ጾ�TѾ��yv,��e?���?��o-�O#���Ӿ����ު)�O����m���4�<P   P   �]�<�B=�ǫ<�s�����b�6�#A������2�.��ra�����rP��T��]bc���0�����-���;�٥���m��P   P   �d��J�<>͎<��G�>&���5�� ��#���G�lc������{��)¿�z��C����J�m|	�ܱ���;�Q���P   P   ����jd.���;:��ŀ�$�f����z��[P��I��ziɿ�K���� �����˿w���H]T�n|	�-���)�P   P   ����Z��\�s�L�
ZN����Г��u��fF������dԿ�	���6t��C���׿x�����J�������P   P   3j�%��Z�R�� ���H�_�ݽ�a��e;L,��͆�ްǿ}	��a)��*7�\�*��C���˿E����0���ӾP   P   `�����@��v�y	���[��gJٽD]9��͢���	�|?]�XS��7�y]��M6��*7�9t�$����z��bbc�S#�P   P   ��پG����@����x�������:��f���Ҿ1(�돁�����o� �z]��a)�!����.¿X���o-�P   P   '��8]��Y����󇾑h��)���Uڅ�jЈ� ��������%:��Ȉ�����:�	��	��K���{��wP����?�P   P   ���-ižo���P�ľ��<���a羡¾oj���^���{��%:�폁�[S���ǿ�dԿ�iɿ���Â���e?�P   P   �4���ž�Y���X�I` ��*B�� B�����ml���^������1(��?]��͆������I��rc���ra��v,�P   P   �fؾ9s��������F�2���t�8��ݜt���2���qj��#����Ҿ��	�R,�nF��[P���G�;�.���P   P   *���"��'k��z4þs���
t��w������ޜt����¾mЈ��f���͢��e;����z�*�������TѾP   P   $,g�Ǵ>���>�Ւ��#�澵A�j����w��:��� B��a�Yڅ���:�L]9��a�ד��o���� ��-A���ጾP   P   �g�+���޽��C	��yJ���A��
t���t��*B�<��,������rJٽm�ݽ��($��5�q�6��v&�P   P   ֩���xW�g�P�1;�����C	��$��t��I�2�L` ��辔h��|���[����H�!ZN��ŀ�Q&������.N��P   P   � W��D)�g�`��(�,;����Ԓ��y4þ�쾂X�R�ľ�󇾸��|	��� ���L����G�;t��x��P   P   ��<r@�<T�;B�`�T�P���޽��>�#k�������Y��n���X�����@��v�Y�R��\����;&͎<�ǫ<��<P   P   L2!=��=�@�<RD)��xW�彺�>��"��2s���ž(iž4]��G����@����Z�kd.��J�<�B=�^!=P   P   �N�=�W�=��I=�x�<�를qy��z	��m�8f��Ǟ��I&ɾ�_��堠��|p�l�����,���<�<5MH=<�=P   P   =�=�r�=�~M=���<����'ý<9��-�� �¾���CV����v(𾨣ľW��5<�6
Ƚ�)���-�<�7K=P   P   6MH=./q=i�J=��<V� �_۽�iT��Ψ����մ�,0��Y9���0����Ӏ�l����X����+�	��-�<P   P   �<�<�Q;=E'==Z�<qF�I�ٽ/Q^�F��0,��m4�-�[�x�s�`Ct��i]�sn6�n.	�$�����c�����)��P   P   �,���f�<)4=Wھ<蘙��V��rR�ta�����i�D�N/|�hc��/˛��.����~���G�u�%�����X�:
ȽP   P   ����h��i<�?v<I]�<3��C�5�*Φ�_,�	)D�!ă�<N��	X��赿����-�����G�o.	�l��5<�P   P   l�G��Y�AKq�	hټ߉�g��wW���1꾃�2��az������w����ɿܺ��������~�vn6�׀�Z��P   P   �|p����6̽De��q(��8iŽ&����g�-�����6�X��ґ��
��� ɿ��ɿ赿�.��j]������ľP   P   頠���i��|O��U��D\�spS�ΒJ��Wb�@H��<�r,���o�����
���w��X��2˛�fCt���0�}(�P   P   �_��*���Q���˾eY���[�ɾ#L��h���y��� ��5���o��ґ�����@N��lc���s��Y9����P   P   O&ɾ����N�ܾ�U�AU�&�m��T��X�iپ�0��5Xþ� �r,�:�X��az�%ă�U/|�5�[�30�HV�P   P   Ξ��29��(�[lF�+����KĿLĿ���s�E�2rﾒ0��y��@龪���2�)D�q�D��m4�ܴ����P   P   @f��%蛾�6۾��E�~���,��q��U��t�E�iپj���DH��2����1�d,����6,����
�¾P   P   �m�VHg�lq��P������Na���$�C�$�q������X�'L���Wb�ŵg�}W��2Φ�}a��P���Ψ��-��P   P   �	����6L���Ⱦ=�R���¿���$�-��LĿ�T�`�ɾՒJ�-��p��N�5�#rR�?Q^��iT�J9�P   P   �y��� ���ȽR����w�j���¿Qa�����KĿ,�m����zpS�CiŽ߉�K3���V��`�ٽv۽�'ýP   P   �를�Dx��.�1)�� �X����?�R�������/���GU�lY��D\�z(��*hټ�]�����F�w� �;��P   P   }x�<}��<�i<�	q�.)��R���ȾR����E�`lF��U��˾�U�Ke��hKq�^?v<8ھ<4�<��<V��<P   P   ��I=';=�u=�i<�.⼉Ƚ�6L�kq���6۾*�Q�ܾ�Q���|O��6̽^� i<"4=:'==]�J=�~M=P   P   �W�=ѻp=';=���<cDx�� ����MHg�!蛾/9������(����i�}��D���h���f�<�Q;=(/q=�r�=P   P   �2�=,��=(/�=�X=�|�<��ټ�װ�\��ͭf�����-��T��a�h�K"�}ⴽD�ql�<��V=bė=b�=P   P   b�=&��=���=�bT=�}<�����ȽN�.�U�y�>L������{ ��KF���W|�;O1���ͽ���aZj<�\Q=��=P   P   cė=k��=hØ=�[U=��Z<��-�+�VM�-۔�2����ݾX�!�޾���-���T�P��-�7�0�@<�\Q=P   P   ��V=���=�a�=I.[=ڹ�<R�+������9a��6��2��N ���R��$	����+�����e�S ��7�ZZj<P   P   ll�<�^P=ݭ{=�vT=#�<$���?轝2`�I���܌��.���1��0:�3^2���k���^˳���e��-񽟩�P   P   N�6	�<F�=MO=u��<�8ʼ�ý�3J��䧾G���)!��A�I�S��FT���B�)#�l���,���W�P���ͽP   P   �ⴽ��N$X����\�>�O���)����*�K���F߾���E�@���\�6g���]���B������0���?O1�P   P   N"��A�˪ӽؽ�.ֽ��ͽ�������s��»��N���/��xR���f�6g��FT�5^2�'	�����W|�P   P   d�h��U�( y��̗�����ѵ���t���O��,a�c����$پ�F��7��xR��\�L�S��0:�U��&�޾OF��P   P   T�� }��s�׾L��o�@��@����վ�%�����w������F���/�H�@��A��1���_龀 ��P   P   �-���񸾝Y���|�d͵��Xο�����*|��3������%��x���$پ�N����-!�2��R ���ݾĢ��P   P   ����X��P�'�S"���H��[.��k.��f��-���+'��������e����»�L߾O������:��	2��DL��P   P   ֭f�����6�*���	��<Xc��.����c�,8��-���3��%���,a���s�P����䧾Q����6��5۔�c�y�P   P   e���RR�~�Ծ�z�_�8�b��f��������c��f��*|��վ��O�����*��3J��2`�:a�dM�Z�.�P   P   �װ��佋�s�����b���,�C����f���.���k.��������t���ཿ)��+�ý @�ӂ��1+���ȽP   P   ��ټ��}Qͽ^d���i=���˿�,�;�b�@Xc��[.��Xο �@�ֵ����ͽd��9ʼB��t�+���-����P   P   �|�<���<�NA�R�ѽ`0���i=��b��_����H�j͵�v�@������.ֽ��>�S��<��<���<n�Z<��}<P   P   ��X==Q=��=���Q�ѽ^d������z�.���X"����|�Q���̗�ؽu���BO=�vT=:.[=�[U=�bT=P   P   $/�=^��=�}z=��=�NA�xQͽ��s���Ծ�6�T�'��Y�y�׾/ y�Ӫӽi$X�A�=׭{=�a�=cØ=}��=P   P   *��=�J�=`��==Q=���<��
���RR�����X����}���U��A���7	�<�^P=���=i��=$��=P   P   �u�=���=M��=�e�=:�X=�bs<3v�y�ʽZ[(�>�]�B�r�_��*���Ͻز��g`<;V=ޠ=χ�=��=P   P   ��=V��=�&�=���=��U=.�x<ި�d(��4���?���[�v8\�iA��������X�e<�R=É�=���=P   P   Ї�=�=">�=��=�gQ=�^8<�c"���ɽk�#�+�[�7ǁ�G#��:Z����]���%�K�ν�_*�r<��L=É�=P   P   ޠ=�M�=�ʼ=�y�=�1X=�?<�
2�ҷ�D;�xH�������ԭ��3���Ȟ�q���u>����Og<�l<�R=P   P   :V=��=3Ҧ=�m�=�>\=��<��A�)ED�W\��hq����;#�׾:�ξ����`��uH���罔_*� e<P   P   �g`<�**=��]=��_=P:0=IV�<p���0�Ž�{9�Cό�����<���^f����&]���`��u>�O�ν�X�P   P   ڲ��sZ��Ğ��;H�i���1���ء���b �t�\4���Y߾F���*������ᾴ��s�����%����P   P   ��Ͻ�]Ž��콑H
�q	�h��ܽ���Ž���QW�9���	̾ k����*�`f��<�ξ�Ȟ���]����P   P   �*���Q��q��Qn˾��jʾݦ��t�L���$�O�:���}������Aվ"k�H���?���&�׾�3��=Z��mA�P   P   _�;J���U
�OyX�����퉿2�W��B	�ѵ���Y��U�Յ�����	̾�Y߾ྭ�;�ԭ�K#��{8\�P   P   C�r��(Ⱦ�-F�⎴����΀����W���eE���ž�3m��U���}�<���`4�����mq������;ǁ��[�P   P   A�]��\Ǿ��^����QE��ր����(oE��(�z�^���ž�Y�S�:��QW�t�Hό�\\��}H��5�[���?�P   P   ^[(��a���D�7��j�`�sZ������¸���a��(��eE�ӵ����$����b ��{9�4ED�D;�u�#�=��P   P   ��ʽ�M����^����C�&��K���?���ø��*oE��W���B	�{�L���Ž塩�@�Ž�A�����ɽt(��P   P   Jv��Ӿ��ړ�bVT���Y����K������������8�W�⦕�'ܽ�������*��
2�d"����P   P   �bs<��;����=ƾGH��`I��Y�(��uZ���ր�Ҁ��퉿jʾw���1�#V�<��<_?<:^8<˄x<P   P   *�X=�-=h�<�kr��ݾHH����C�o�`�WE���������q	�i�B:0=�>\=�1X=�gQ=~�U=P   P   �e�=wG�=v�_=����kr�=ƾeVT��^��>�����鎴�XyX�[n˾�H
�z<H���_=�m�=�y�=��=���=P   P   J��=7�=T�=z�_=�<���㽱ړ����D��^��-F��U
��q��ɋ�.Ş���]=0Ҧ=�ʼ=>�=�&�=P   P   ��=˹�=9�={G�=�-=q�;��Ӿ��M��a���\Ǿ )Ⱦ@J����Q��]Ž�sZ��**=��=�M�=�=T��=P   P   �a�=�W�=�A�=��=8��=K�:=�^b8�%n�w<��1�DkF�!�2�����@w��ͺձ6=��=P��=HN�=�s�=P   P   �s�=)z�=���=�/�=}�=1�X=k��<���� �����ս�������׽<ǋ���̼�ˈ<W�U=��=���=���=P   P   IN�=.�=H��=W��=ѣ=�KV=\�<�ü�(��,`Խvf�Lw��*�X�ֽ�P��T�ϼH�<�4R=|k�=���=P   P   P��=,b�=���=���=5ؤ=�W=�y<+��	 ���@���Q!�J�5���5��"�����"��R7 �[3^<�4R=��=P   P   ��=�d�=���=ޑ�=V��=�O\=kݐ<y�켐3��X��:��Z�(�f���[��|<�����y��T7 �C�<U�U=P   P   ձ6=mt=���=�w�=��x=�H>=�"�<D�����^
��C���p�Z���|���wr��yF����$��\�ϼ�ˈ<P   P   ��ͺ+1�;M_�9���C�:�M�;׆�:&s��~���K����8���o����G���!a���wr��|<������P����̼P   P   �@w�'��������/ �}m�u���ܑ���Oh��n��O3ν�W�{nX�Z���f%��H���}����[��"�]�ֽ>ǋ�P   P   ����hN��5����T.�o#ﾖ���>vJ�@/����ν@���1�@�c�Z������\���-�f��5��*���׽P   P   �2�3j��{o��8���Ӧ�粦�〿*���`���$.�6���V��1�}nX���o���p��Z�O�5�Pw���P   P   AkF�S�ҾC�f��SٿC� ���7�w� �Dٿ�uf�e*Ѿ��B�8���B���W���8�%�C��:��Q!�{f����P   P   1��Ѿ/e��Q����n�JY���s��!\o�� �E���f*Ѿ�$.�ŠνW3νV���^
�_��@��9`Խ��սP   P   z<��0/����d���jه�?����W��'��R���� ��uf��`��H/���n�����������3�� ���(��*���P   P   �%n�ƛI����x�ֿYm��j��П������'��$\o�Dٿ-��EvJ��Oh�Js��o�����_��7�ü���P   P   �#b8h�� ֥�s6}�؋�x���C���џ���W���s��{� �〿����瑤����:�"�<Bݐ<��y<�[�<B��<P   P   =�:=b>�;x��P�龮C���4�y����j��A���MY����7���x#ﾄ���SM�;�H>=uO\=m�W=�KV= �X=P   P   2��=��w=�58;�"�����C��ً�^m�mه���n�I� ��Ӧ�Z.��m�	
�:��x=P��=.ؤ=ѣ=w�=P   P    ��=�ƺ=3�=��w9�"�R��w6}�|�ֿ��V���Sٿ�8����/ �E����w�=ڑ�=���=R��=�/�=P   P   �A�=��=5��=5�=.68;�x��"֥������d�4e��L�f��o��5������X�9���=���=���=E��=���=P   P   �W�=���=��=�ƺ=��w=�>�;h��țI�4/���Ѿ[�Ҿ9j���hN�1����0�;it=�d�=*b�=.�=(z�=P   P   y� >	��=�=��=��='�=���<�%Ἒڰ��h
�^������o��t(�9��<ht�=l�=l��=kH�=?��=P   P   @��=m��=���=Һ�=J��=
s�=�@S=v��<?4����A�If��-��b�E��	��;��<�O=Xe�=��=e��=M��=P   P   kH�=���=���=��=#2�=�S�=�9d=%m�<b=1�(l�\G�3�d��uI�Hg��Ou����<f�`=v�=�U�=e��=P   P   m��=�Z�=��=�W�=W�=�Ӥ=4Zd=��<�{��G����o��w��o���r�^�xd޻c��<v�_=v�=��=P   P   l�=�/�=8��=��=�={á=��f=��<! �d>-��I���R���(˽��������QZ3��*�a��<e�`=Xe�=P   P   it�=�&�=i��=v,�=�=�_�==W=�;�<�ș�+�b坽Vֽ�\���-����ؽ/O��RZ3��d޻���<�O=P   P   D��<�<�B�;Q�:lX�;��<�P�<�ץ<��(�
�����-ս���
������ؽ����c�AOu�;��<P   P   `(�C��Z��������5�+��%|ڼtl��z༦�g�����(�� 
��
��-�������r�Rg���	��P   P   �o����<�����������ﾺI��;�9�rm��8�gA<��[���ƽ�(���\���(˽t���uI�a�E�P   P   ���}Ý�����+�������⦿�怿|"�)$���n�GE�� �W��[������-սVֽ�R���w��=�d�-��P   P   Y��|~Ⱦ��d�K�ؿ1f �7�rr �ݭؿ@�d��qǾP��IE��lA<���g����j坽�I���o��\G�Jf��P   P   �h
��Ǿ�>����W�m�������5n���۲���qǾ�n�8��z�6�
�,+�w>-�Y��Gl��A�P   P   �ڰ�)�����b��{����A����|���U���܇���C�d�+$��xm���l�z���}ə�X! ��|��p>1�V4��P   P   �%�}�7�'��տ]�k���������� V���5n��ؿ"�A�9�C|ڼ�ץ<�;�<��<���<m�<[��<P   P   ���<�����2���}�f��5����������|����ur ��怿�I���+���P�<�<W=��f=$Zd=�9d=�@S=P   P   �&�=�:�<����V��G&4��5������C������7��⦿����5��<�_�=uá=�Ӥ=�S�=s�=P   P   ��=��=n�<qu��p��V��h�a�k����^�m�7f ���������W�;�=��=W�=2�=E��=P   P   ��=({�=��=F��;ru����}�$�տ�{���S�ؿ�+����� ���N�:r,�=��=�W�=��=Ϻ�=P   P   �="�=_i�=��=s�< ��2��+���b��>����d��������k��B�;e��=6��=��=���=���=P   P   ��=��=#�=*{�=��=�:�<������7�-����Ǿ�~Ⱦ�Ý���<� C��ڕ�<�&�=/�=�Z�=���=l��=P   P   �P>�1>:��=j	�=�`�=���=֏-='���b��8ȽTP�c�ʽȪj��2��}�(==H�=B��=�%�=��=�I>P   P   �I>bG>���=���=�U�=�J�=Hk�=�9=��<�e�ۑɼ`A̼�p��׀<�$6=�.�=�=��=��=��=P   P   ��=<��=�?�=��=q%�=D��=ǐ�=3�o=��=�Ǌ<�k0;Ͻ,���;�؅<��=�m=u��=���=���=��=P   P   �%�=�_�=Ȓ�=��=�='�=�,�=��w=�� =��<�^Y;{[������:;�~�<��=��t=���=���=��=P   P   B��=���=-R�=�2�=@�=f�=��=�y=�1=V2�<(G(����ۑ������W�m�<��=��t=u��=�=P   P   >H�=���=���=b5�=*�=���=/�=�,s=,�#=D��<���C���^(�d�L���jϻm�<��=�m=�.�=P   P   ��(=�Z�<Ccw<nE<cс<�~�<k�/=�>=�=Au�<�0�SF����0-��}�O����W��~�<��=�$6=P   P   �2�� D�y�ȽQ���G�'Ž��;�,�`��}�<���<���;�.l����l�+�2-�h����[�:;�؅<؀<P   P   ��j�g��V򎾺�;c4�,�̾�Ѝ��$�E_���xL�;�i�4��������d(�葦����n�;�p�P   P   Y�ʽ0����d��Y��A��B.��ؤX�����a��	"Žd^���Ǐ�%�i��.l�aF��T���ֺ��[���,�ZA̼P   P   KP�
��sA@�_P���:���5I�%g��@��3��i��h^��XL�;{��;�1�X����G(�^Y;-k0;ّɼP   P   �8Ƚ�=��uX��#�]�B��}�;~�s"C�
��>Y��3��"ŽK��湘<.u�<.��<>2�<��<�Ǌ<�e�P   P   �b�~́�с>��"濮!]����-b����Rt^�
迁@��a��E_��}�<�=!�#=�1=�� =��=��<P   P   '�����(�y��� A�����{����1����u"C�(g������$���`��>={,s=�y=��w=(�o=ۨ9=P   P   я-=�z7�i+����T��=�\{����{���.b��@~�8I�ޤX��Ѝ���;�a�/=*�=���=�,�=�=Dk�=P   P   ���=G��<9��$ȾkG���:�
\{���������}���F.��3�̾3Ž}~�<���=f�=#�=@��=�J�=P   P   �`�=x�=/�<�a���lG���=�� A��!]�b�B��:��A��m4��G�Eс<*�=@�=�=m%�=�U�=P   P   h	�=[��=�
�=R�:<�a�&Ⱦ��T�}���"濦#�fP���Y�Ù;Z��,E<^5�=�2�=��=��=���=P   P   9��=:�=I1�=�
�=/�<
9��l+��,�ׁ>�uX�{A@��d�]򎾉�Ƚcw<���=+R�=ƒ�=�?�=���=P   P   �1>;!�=:�=]��=z�=J��<�z7�����́��=��
��6���p��D��Z�<���=���=�_�=;��=aG>P   P   �f�=�k�=��=��=e �=K[�=:Q=�}I<���낽����߄��)��h�3<�=M=r�=K��=���=�f�=Ƣ�=P   P   Ǣ�=��=X��=���=��=��=��=%�p=�=�/r<��;��:Oih<��=?@n=�Ϣ=�u�=���=��=��=P   P   �f�=z�=�x�=2��=i��=m��=�o�=�=h�m=+�/=h<=��<�G=e-.=�k=�	�=�Ƶ=j	�=D��=��=P   P   ���=��=�.�=S�=���=���=���=>�=_q�=��K=�=t=��=�:=GJ=�]�= ޞ==j	�=���=P   P   L��=1a�=Pe�=w��=���=w��=�]�=G�={w�=$�M=^�=p��<8��<e��<�=�!K=��= ޞ=�Ƶ=�u�=P   P   r�=���=�0�=��=W�=8a�=�=�s�=�=y/O=w	=)}�<�'�<��<�~�<��=�!K=�]�=�	�=�Ϣ=P   P   �=M=T�=��<��<ep�<��=1GS=�t=�)r=&�O=�=#�<�+�<ˬZ<���<�~�<�=EJ=�k=B@n=P   P   ��3<r�8�����ɽJ�Ƚ�錽͗Ҽ=�T<I =��5=��#=޼�<\��<�$_<ƬZ<��<`��<�:=e-.=��=P   P   �)����བ�X�vl��󧮾�ؚ�ۈV�f�۽�t�<��<�x
=GK=m�<Y��<�+�<�'�</��<��=�G=bih<P   P   ߄�o�E� Ǿ���6�H�A�H��F�h�ž�C�������;8��<FK=ؼ�<#�<}�<d��<o={��<���:P   P   {���Ů|����~� N��ѿ�X����~�����z�����;�x
=��#=�=q	=V�=��=d<=�;P   P   �낽��{�m������-��{-���-��~��~���|��z����3��<��5=�O=r/O=�M=|�K=&�/=�/r<P   P   ����B�b���P��|��%`�k����`����~������C��t�C =�)r==ww�=[q�=b�m=�=P   P   �}I<�Uڽ��þ�{�)0�	K_������ڑ���`��~���~�k�žn�۽�T<	�t=}s�=C�=:�=�= �p=P   P   8Q=��μ�S����������+��~�����n����-��X���F��V��Ҽ(GS=�=�]�=���=�o�=��=P   P   J[�=
B=ڸ��#����E���Ϳ��+�K_�)`��{-�ѿG�H��ؚ��錽|�=4a�=t��=���=j��=��=P   P   c �=à=N�<G��������E�����+0�����-�N��=�H�����W�ȽLp�<S�=���=���=g��=��=P   P   ��=�]�==�=Bؚ<H���$�������{��P��������~����}l���ɽ��<���=u��=S�=1��=���=P   P   ��=ǘ�=�$�==�=N�<ܸ���S���þf��r�� Ǿ��X�D�����<�0�=Ne�=�.�=�x�=W��=P   P   �k�=�
�=ǘ�=�]�=à=B=��μ�Uڽ�B���{�Ю|�y�E���:r�J�=���=0a�=��=z�=��=P   P   H�=�E�=�_�=�K�=P|�=I�=$:S=�&�<�f��o'��R���)�WLu��<��P=���=x��=	��=0��=�{�=P   P   �{�=6p�=9�="�=Ѓ�=���=R��=��{=R�-=�C�<�|<�Tz<S��<��+=/Dz=��=�~�=���=�6�=�X�=P   P   1��=��=���=�R�=H�=��=�g�=�0�=́�=G[=:�7=��*=�)7=��Y=��=���=���=���=���=�6�=P   P   
��=��=���=��=��=uF�=j��=���=;4�=}�=�a=��N=$mN=%�`=go�=Oi�=E��=�ֺ=���=���=P   P   y��=`��=���=�h�=�l�='��=VF�=+K�=q�=f.�=j=�9R=�vI=�}Q=ߗh=U)�=��=E��=���=�~�=P   P   ���=#�=�/�=坏=T�=;�=��=H��=�U�=���=zUk=�zN=�>=�==��L=��h=U)�=Oi�=���=��=P   P   ��P=��=I�<Ag�<���<	�=�SV=}	�=:��=�ւ=Z{l=ߑO=�c9=D�0=�8=��L=ߗh=go�=��=2Dz=P   P   �<�0i���E�!���3����@��dM��'�<VV3=�`=U-f=��U=�@=�1=C�0=�==�}Q=$�`=��Y=��+=P   P   +Lu�NR�����R2a�q|��`�g��筚��O��%�<��>=�)T=5xM=�@=�c9=�>=�vI=#mN=�)7=\��<P   P   ��)�SP�����ܾ{��غ���۾�Ս���� �"َ<62=�)T=��U=ܑO=�zN=�9R=��N=��*=�Tz<P   P   ��R��7�ۀƾī*��o�����n�=*�Ifžq=5��I� َ<��>=R-f=V{l=vUk=j=�a=8�7=�|<P   P   zo'��6��wܾ|�T��Ш��׿�׿ᨿw�T���۾r=5�� ��%�<�`=�ւ=���=c.�={�=D[=�C�<P   P   �f�	���6ž�8T�=���B�	�=C���	��A��x�T�Jfž���O�QV3=8��=�U�=n�=84�=ˁ�=Q�-=P   P   �&�<�s���5��)��ا�'4	��d1���1���	�ᨿ=*��Ս����'�<{	�=E��=)K�=���=�0�=��{=P   P   #:S=��P���/�پ��l��zտƪ��d1�?C��׿��n���۾l���dM��SV=��=SF�=h��=�g�=Q��=P   P   H�=� =Ϡ=��\���������zտ(4	�D�	��׿��ۺ��`���@��=;�=%��=sF�=��=���=P   P   O|�=�`�=Wt�<k���R�w������l��ا�A����Ш��o���z|��3�����<Q�=�l�=��=F�=΃�=P   P   �K�=���=��=n��<l����\�1�پ)��8T���T�ɫ*��ܾ[2a�+��+g�<❏=�h�=��=�R�=!�=P   P   �_�=Y<�=�P�=��=Vt�<Ҡ=�����5���6ž�wܾ�ƾ��������E�5�<�/�=���=���=���=9�=P   P   �E�=-��=Y<�=���=�`�=� =��P��s����"�6��7�ZP�XR���0i���= �=_��=~��=��=5p�=P   P   �n�= ��=���=�%�=F�=�ԇ=�/5=�	�<vM8� ��*��z	��A�m��<��3=`��=��=�}�=S:�=��=P   P   ��=>��=p�=���=6�=컨=� �=��b=� =#C�<���<-��<u>�<�==��a=0؏=�=��=S�=�=�=P   P   T:�=�E�=<I�=x:�=�.�=b�=��=t�=8~=~�V=&:=�/=z9=�V=DW}=Wy�=�7�=�״=� �=T�=P   P   �}�=cq�=��=hռ=ș�=?p�=Թ�=%�=+ۑ=U�=n�l=Z�^=�^=�Al=sk�=�<�=�ӟ=��=�״=��=P   P   ��=r�=�ޥ=!�=�=Ω=k�=�="ݖ=��=�
=��n=�h=�n=��}=w�=�ڕ=�ӟ=�7�=�=P   P   a��=e?|=�!p=w�p=Q�~=F�=���=TV�=���=ۄ�=?�=��r=�7h=%�g=39q=>�=w�=�<�=Wy�=1؏=P   P   ��3=n�<]�<�<jʦ<m�=H9=�gg=�4�=���=���=��s=J�g=ːb=(bf=39q=�}=sk�=FW}=��a=P   P   z��<p8N��(�Mq�(o���"���1�O"�<�}&=pW\=1Pq=�q=j=Ic=ʐb=$�g=�n=�Al=�V=�==P   P   �A� ����Y��N3��MG��1�����}�1��4�<��@=^�c=Fl=j=I�g=�7h=�h=�^=z9=|>�<P   P   �z	�H轮�a�����ϾtQϾ%����N^�b��B���Ɨ<`26=]�c=�q=��s=��r=��n=Y�^=�/=5��<P   P   �*�3��#��;�����.�!BB�K.������*��XB�����Ɨ<��@=/Pq=���==�=�
=k�l=%:=���<P   P   �1=����%T�os��Ϛ��{��>#r�l�a���XB�G���4�<nW\=���=ل�=��=S�=|�V=%C�<P   P   gM8�xu�u���/�f����1ȿ���7zǿ!6��l��*��e��B��}&=�4�=���= ݖ=)ۑ=8~=� =P   P   �	�<m���t�_�i�����r�;0ȿ������8zǿ?#r������N^�}�D"�<�gg=RV�=�=#�=r�=��b=P   P   �/5=��A��W��ʽ��.�����J�������俼{��M.�(���������1�H9=���=k�=ҹ�=��=� �=P   P   �ԇ=s	�<Z\$�!�1���ξ��A�����<0ȿ�1ȿ�Ϛ�$BB�xQϾ�1���"�g�=F�=�ͩ=>p�=a�=뻨=P   P   F�=O|=J�<�m�F���ξ.���r�h���os���.���Ͼ�MG�*(o�[ʦ<L�~=�=Ǚ�=�.�=5�=P   P   �%�=��=�o=���<�m�"�1�̽��l���1�(T�A�����!N3�[q���<r�p=�=gռ=w:�=���=P   P   ���=��=7�=�o=J�<]\$��W��w�_�x������#����a��Y���(�M�<�!p=�ޥ=��=<I�=o�=P   P    ��=���=��=��=O|=r	�<��A�p���~u�5=�7��H�����8N�a�<a?|=r�=bq�=�E�=>��=P   P   �,�=|1�=q+�=�a�=�U�=�uQ=���<�J�;K����=#�PB�/�#�������;���<��Q=���=ڻ�=�|�=�^�=P   P   �^�=6W�=ʿ�=W �=���=���=��g=p�/=�9�<��y<���;bu�;�Nw<6��<�/=[�g=�=�ʚ=�!�=&֪=P   P   �|�=��=���=.E�=Am�=7�=�܋=X�w=��S=}Q1=�R=[�=�=��0=�S=P3w=���=!��=G@�=�!�=P   P   ڻ�=kǛ=��=��=�I�=���=P�=��=�M~=l#g=~}S=HH=��G=�R=a@f=�5}=�~�=�G�=!��=�ʚ=P   P   ���=;��=g��=��=�y�=寋=b��=���=�A�=��{=o�l=~a=a�\=��`=��k=�Qz=$C�=�~�=���=���=P   P   ��Q=��;=�m.=�;/=E>=)�T=8Ek=d�z=W<�=}=Kt=��j=�[d= �c=`i=�r=�Qz=�5}=Q3w=]�g=P   P   ���<9�<�&�;x�*;HZ�;�Փ<Z�=�4=pX=�dj=�n=��k=Uf=��c=�se=`i=��k=a@f=�S=�/=P   P   ��;b\���BG�����u�����A�82��9|�;�w�<A�6=,�W=\ad=�f=��d=��c= �c=��`=�R=��0=<��<P   P   u���������ض,��c>��+�����R�������Y�<�=HM=�G`=�f=Tf=�[d=a�\=��G=�=�Nw<P   P   (�#�,���dV�� ������T���$��0R���߽ņ�B#!<�	=GM=[ad=��k=��j=~a=GH=\�=|u�;P   P   �OB���ܐ���|P&���:�f�$��i쾆獾Y��^Z5�?#!<�=*�W=�n=It=m�l=}}S=�R=���;P   P   �=#�p��8��/�IRs�����<��$6p�Z���ʜ�Y��ǆ��Y�<?�6=�dj=}=��{=k#g=|Q1=��y<P   P   D������*����D�����޿] ��ܿ#k��[���獾��߽�����w�<mX=V<�=�A�=�M~=��S=�9�<P   P   �J�;3G����U�V���s��G߿O&�IP%��ܿ&6p��i�2R�"R��|�;�4=a�z=���=��=V�w=o�/=P   P   ���<����4�������&�����X� O&�^ ��<��h�$��$�����C2��W�=5Ek=a��=O�=�܋=��g=P   P   �uQ=w'�<k�F���,��t¾�b<�����G߿��޿�����:�W���+���A��Փ<&�T=䯋=���=7�=���=P   P   �U�=;=[-�;51���9?��t¾��&�
�s�E���MRs�P&������c>�y���Z�;A>=�y�=�I�=@m�=���=P   P   �a�=��=O-=�(;61����,����Y���1���� ��ܶ,������*;�;/=��=��=-E�=W �=P   P   p+�=�>�=�ǂ=O-=W-�;m�F�4����U�,���;���ܐ��dV�%����BG��&�;�m.=f��=��=���=ɿ�=P   P   |1�=���=�>�=��=;=v'�<����5G�����s���2�����q\��.�<��;=:��=jǛ=��=6W�=P   P   5�=��=줂=(�l=�mD=��=�V<0C6�����_�V�}�A4`�:p��7�M7V<�9=�E=��m=h��=�,�=P   P   �,�=�(�=J��=��=�m=�*N=r�"=���<��L<���9���:n���D9�NK<u�<f�"=�+N=6�m=���=���=P   P   h��=�p�=���=�$�=�-z=B�k=�{U=t�8=
�=^�<���<ձ<�U�<���<9)=�8=i�T=U"k=3�y=���=P   P   ��m=W�l=m=gan=,�n=sfl=V�d=E�W=�IF=�T3=�#=�P=�=J�"=Ǎ2=�,E=Y�V=��c=U"k=7�m=P   P   �E=�`==,�:=CO>=#�F=GaP=�CW=�X=J�T=��K=ыA=�l9=*6=v�8=B�@=�1J=�R=Z�V=j�T=�+N=P   P   �9=wT�<)��<�4�<��<5�=�C&=ͫ;=�^H=��L=��J=̆F=URC=�B=/eE=��H=�1J=�,E=�8=h�"=P   P   Z7V<��W�l<��){�fm1��o�9�>l<7�<l#="�6=��C=kzG==cG=��F=\SF=/eE=B�@=Ǎ2=:)=z�<P   P   �7�[u��鄽qn��?D���災�r���?�h<g�<EW'=�C<=��D=�?G=��F=�B=v�8=J�"=���<�NK<P   P   5p�%�9��!;�V�L��=9��>
������7�]�;v6�<�2=�j9=��D==cG=TRC=*6=�=�U�<�D9P   P   ;4`�����d�"���K7̾ ?˾#B���_�Hq����R�R���A�<�2=�C<=jzG=ˆF=�l9=�P=ձ<"n�P   P   Q�}�!��혾����w6���N��4�����9������so�V���t6�<DW'=��C=��J=ЋA=�#=���<���P   P   ��_���c֨��<!�!k���࿿|�����K�����������R�G�;g�<!�6=��L=��K=�T3=^�<v��9P   P   ��k����k!�l��;���=6�����ꞿK���9��Iq���7�7�h<k#=�^H=I�T=�IF=
�=��L<P   P   *C6��㫽G e�sR�����od�6�i�3h����������_�������2�<˫;=�X=D�W=s�8=���<P   P   �V<B����o<��oY7�L ¿�e8�7�i��=6�}����4�$B���>
��r��>l<�C&=�CW=U�d=�{U=q�"=P   P   ��=Y��ҩ��2<���;UtQ�L ¿pd�<���࿿��N�?˾�=9��災�m�93�=EaP=rfl=@�k=�*N=P   P   �mD=�,�<E�B��'����N���;pY7����l��#k��z6�N7̾Y�L�BD��xm1����<!�F=+�n=�-z=�m=P   P   (�l=|6<=tԿ<黃��'��2<�p<��uR���k!��<!�����$����!;�un���){��4�<AO>=fan=�$�=��=P   P   줂=��k=m�8=tԿ<G�B�ө����I e���e֨��혾��d�9��鄽�<�#��<*�:=m=���=J��=P   P   ��=G�=��k=|6<=�,�<%Y��D���㫽l���!���*�au���W�rT�<�`==U�l=�p�=�(�=P   P   �K=-G=��9=մ =�S�<!p<k�����o1U����M�����PU���缀Ɵ��r<�r�<�R!=�J:=�qG=P   P   �qG=�mG=I`B=��6=ٷ"=��=}�<4�<6/���s������Ż��郼cS���<<@�<��=3�"=��6=lB=P   P   �J:=m;=�r:=�57=�/=s="=Y�=��<��<��]<q@<l��;)<C6\<��<%��<zE=�!=]-/=��6=P   P   �R!=z ={e =�"=��#=��"=_�=$�=x=��<���<���<u+�<���<�P�<�_=��=�=�!=4�"=P   P   �r�<���<��<;��<n��<$=%�=��=`{=��=�<	=Lq=�1=^�=�#=BY=�=��={E=��=P   P   �r<��<O�;��;�2<3<Q{�<���<2�=��=�="B=��=�c=�)=�(=BY=�_='��<?@�<P   P   jƟ������O�)!	�d������ֱg��)<���<g[�<�)=� =�A=K�=O7=�)=�#=�P�<��<�<P   P   ���?e��צ���ƽ�lŽ�Σ��]��׼D(+��zt<1/�<^1=�T=�"=K�=�c=^�=���<H6\<QS��P   P   PU��˽���y�H�>�Y��F����SXŽ�J�Ƹc��k"<3��<;g=�T=�A=��=�1=v+�<.<�郼P   P   ��������p�D�����о�Ͼ�=����k���vG���ȧ��M<3��<^1=� ="B=Kq=���<t��;Ż�P   P   M��Ĵ+��,��pt�~�8�=�Q���6�5 ��U��wO&�� ���ȧ��k"<//�<�)=�=�<	=���<t@<����P   P   �����+�签ǲ#�����jĿ� ÿ8������o��xO&�wG��ʸc��zt<e[�<��=��=��<��]<�s��P   P   m1U���_Y����#�������=�Q��١����U�����J�](+����<1�=^{=x=��<//��P   P   ��̽�uq�����G��cG���s�O
r�Q�8��6 ����k�UXŽ�׼�)<���<��=#�=��<5�<P   P   f�����e��d�0���/!:���ƿr=?���s� =�� ÿ��6��=������]���g�N{�<$�=]�=X�=}�<P   P   !p<�ĝ�� ��z�I��Ҿa�T���ƿdG�����jĿ?�Q��Ͼ�F��Σ����+<#=��"=r="=��=P   P   �S�<�<<|�����Ƚ�0\��Ҿ0!:��G����������8���оA�Y��lŽk��2<k��<��#=
�/=ط"=P   P   Դ =a��<�d�;>����Ƚ{�I�1��������#�ɲ#�qt�F���|�H���ƽ-!	���;7��<�"=�57=��6=P   P   ��9=�=���<�d�;}���� ���d��uq�aY��
签�,����p�����צ��O��N�;��<ze =�r:=H`B=P   P   -G=1�:=�=a��<�<<�ĝ���e�̽��»+�ƴ+�����˽Ee�������<���<y =m;=�mG=P   P   �=U�<�w�<��<�I=<��%����o|/�Pj��䭦��������4j���R/�a���w�:?<�a�<�+�<���<P   P   ���<\��<�K�<Ύ�<Ø�<��m<�;ۄ�����A���<�#X����B���f�ﻨ��;�m</{�<3~�<�^�<P   P   �+�<d>�<���<BU�<k��<~ͳ<�	�<��8<�w�;,��s�߻<T�_�E4�^]�;�(6<	��<�s�<v��<4~�<P   P   �a�<���<e(�<C�<���<9�<��<uf�<毅<�zT<^$<�<^<a"<��P<�l�<zњ</9�<�s�<0{�<P   P   =?<��<��<�<)�E<�v<D!�<�-�<ӹ�<���<Tݗ<)��<�)�<֎<���<��<6՟<{њ<
��<�m<P   P   �w������E�}�B�B��Cܺ�|�;ݽC<�<���<���<���<)��<׽�<�^�<K;�<��<�l�<�(6<���;P   P   ]��H~���6��E�sx4��>	�/١��ƻ1#�;�`<�<�D�<���<�i�<h�<�^�<���<��P<f]�;Z��P   P   �R/��ƌ�2��mڽ�ٽk:��8��Ү'�����b"^�J�3<R��<
n�<҃�<�i�<׽�<֎< a"<54�>���P   P   2j���
޽I���G�6�V�O�E���J1ؽ�_~�����'��֒<S�<
n�<���<(��<�)�<_<W����P   P   ����x�g k�����9��$^��ݏ��Xf��d�Y����AG�Ւ<Q��<�D�<���<(��<�<8T�!X�P   P   ������-�-����꾰� �HS4�^
�J��HՒ�l�(��լ����'��H�3<�<���<Tݗ<^$<m�߻�<�P   P   ⭦�I�-�̛���O�ԯk��̜����*h��X�����l�(�Y����鼏"^��`<���<���<�zT<'���A��P   P   Nj��V���Y���y��ۇ��~Ή]
���޿WO���X�HՒ��d��_~�����)#�;���<ҹ�<寅<�w�;���P   P   m|/��k޽%�k�ł��l�4[��.�Ԓ-���޿+h�K��Xf�L1ؽԮ'��ƻٽC<�-�<tf�<��8<ل�P   P   ���hB���k ��i��Y�!��;�����.��]
����_
�ޏ����:��3١��|�;B!�<��<�	�<�;P   P   ��%�Η��;��&I�!�¾��6��;��6[⿠~῍̜�JS4�%^��P�E�m:���>	�(Dܺ�v<8�<}ͳ<��m<P   P   �I=<1Z��#9��Uܽ�*Y�"�¾Y�!��l��ۇ�ׯk��� ��9��8�V��ٽvx4� B�$�E<���<j��<�<P   P   ��<Z�<�jM�QI��Uܽ'I��i��Ƃ��y��O���������G�pڽ�E���B��<B�<AU�<Ύ�<P   P   �w�<V�<C6	<�jM��#9��;���k �'�k��Y��͛���-��j k�K��4����6���E���<c(�<���<�K�<P   P   
U�<�+�<V�<Z�<2Z�ϗ�hB���k޽W��K�-���-��x��
޽�ƌ�K~������<���<c>�<\��<P   P   l�u<��d<�0<ï�;{��m̍�`�J-Z�ν��m䰽[黽^谽/���Z�j)��3��*����ݠ;o1<7e<P   P   7e<_We<КP<�(#<�`�;��Ǻ�-�l���LG�0,��B�nC��[,�0���I��L0.�a�ͺ��;��"<�`P<P   P   p1<rN5<�)2<��$<w	<w��;��:RC��PZ)��惼��(�B����턼&�+�5����N�:�®;��<��"<P   P   �ݠ;��;O��;j�;���;�g�;\?�;�hY;�Yc:�&��pΏ��g������T��b��L,:�DD;�r�;�®;��;P   P   $���%�λ�廕ȻFE���ڌ�65�:|e;S��;B1�;�{;��R;��>;�7J;_5k;C��;﵂;�DD;�N�:N�ͺP   P   �3��x����ռ�DԼ/���v���=K!�V�n���:G1�;��;#&�;E��;�t�;���;�W�;D��;^,:1���I0.�P   P   h)���<�,�a�l�n��}_�I39�V���������+��|Q�;)o�;�<��<�<���;a5k;]��#�+��I��P   P   Z�]g��̫Ľ�*ݽ�Fܽ�H½�/��t\S�����-+u��@h��]w;�< 6<��<�t�;�7J;T���턼/��P   P   .���T�YN�)_8��VD�"�6���۽�2����$��󚼗����i;�<�<D��;��>;����@����[,�P   P   ]谽���&T�u��u񢾞Q��튾�mP�s[�#w����:�� ������]w;'o�;!&�;��R;�g��&�lC�P   P   Y黽S#�����e��������3���$���Ռ��y^�����:��󚼸@h�yQ�;��;�{;oΏ����B�P   P   l䰽�\#�c!����/q)�WhV�kjU��T'�X���;��y^�#w����$�/+u�;��C1�;?1�;�&���惼0,�P   P   ͽ�����48��~�G�>����⛡�pߊ�H�;�X��Ռ��s[��2�����������:O��;tYc:OZ)�KG�P   P   I-Z�pTཊ�T�������)�6|��[��ss��pߊ��T'�%����mP�۽u\S�����a�n�|e;�hY;SC��k���P   P   `��՛����B��������W�����[��㛡�ljU�5���튾���/��X��@K!�"5�:Y?�;��:�-�P   P   l̍���=�P�Ž=|9�(��>�	���W�6|�����YhV����Q��#�6��H½K39�x����ڌ��g�;t��;��ǺP   P   {���`��b�c�A߽�2F�(��������)�I�>�0q)�����v��VD��Fܽ�}_�2���ME�����;~w	<�`�;P   P   ¯�;"ֻ%ټ��q�A߽>|9�B�����������e��u��+_8��*ݽo�n��DԼ�Ȼe�;��$<�(#<P   P   �0<�1�;�q�%ټc�c�P�Ž�����T�58��d!�����(T�ZN�ΫĽ/�a���ռ���J��;�)2<ϚP<P   P   ��d<�@3<�1�;"ֻ�`����=��՛�qT�����\#�S#����V�^g����<�x��,�λ��;qN5<^We<P   P   ����������~��������'�2�}t��ڙ��'���˹��*���ڙ�1|t�g�2��D�!a�����N���P   P   ����Z���š������{�x���9���,���M��g`��z`���M�;'-�x^��s��5*}�����"��#�P   P   L�����x�ڃ����Neӻ�=�]�R�^ɐ��㻼���� ���` �����vM����U�&Z�Sٻ�"��P   P   ��d ���^��}g�"B����32���S�L1y��P��SW���e��ف|�VtX��E7��!�%Z����P   P    a������f���_�������u�y�M�DJ/��U�(�!���$���'���&�_�"�q� �� &��E7���U�3*}�P   P   �D�/�KG�)���c
��4��к�����8N�t,�$��ɻˮ��%,����л����q� �UtX�uM���s��P   P   f�2�k�\��.{��ނ�3ey���Y�(�.��X�����o�o����û�y��t�s�������л^�"�؁|� ��x^�P   P   /|t�3���8���lԽo�ӽ�S��a�����n���'� ܼGL�����B����k�u�s�&,����&��e����9'-�P   P   �ڙ��ֽn&
���!���*�'� ��u�k�ҽ/,��-�G�S	��������B���y��̮����'�SW��_ ���M�P   P   �*��̍���5�<�e���������6�c��@3��� �zͬ�ГY��������ûɻ�$�~���z`�P   P   �˹�<D���X�`����ķ�_�ž���j7���wU��G�N8��ГY�S	��GL���&��"���P���� ��g`�P   P   �'��dI��f��s�����x�	��	�ڟ�w��h�b��G�zͬ�-�G� ܼp�o�u,�)�L1y�����M�P   P   �ڙ�����,Y�����������'���9�j&�����w���wU��� �0,����'�����9N��U���S��㻼��,�P   P   }t���ֽj76�2K��%O�q�'��'Q��P�j&�۟�k7���@3�k�ҽ��n��X�����EJ/��32�^ɐ�9�P   P   '�2�������
���f����
�s�:��'Q���9��	����8�c��u�a���)�.��к�{�M���^�R�x���P   P   ���g]�k½�"�Pɂ��Ǿ��
�r�'���'�y�	�`�ž����(� ��S����Y��4��u�$B��=���{�P   P   ����\���|��ս6�+�Pɂ��&O龖������ŷ�������*�p�ӽ5ey��c
�����~g�Peӻ���P   P   ~��O��S������ս�"���f�3K�������s��a���=�e���!��lԽ�ނ�*��	_��_������š�P   P   ����\"��᧼S���|�l½��
�k76��,Y��f���X���5�o&
��8���.{�LG�g�����ڃ�]��P   P   ���(�\"��O��\���g]�������ֽ���eI�=D�͍��ֽ3��m�\�0�����f ���x�����P   P   =^V���e�������������O��Ɓ��Q��O4���Ų�7���\��9ȁ�O�u����Lc�����pe�P   P   pe��!e���x�A��d^����ܼ{]
��I*�t�I��d��s��*s��@d�P>J��*�ڽ
�K�ݼ������jay�P   P   �����������ӏ�]&��Jׯ���ʼI*켏O�z����$��*)��$��[����%��m̼�`����������P   P   Lc������(��j�����e���K��"����xɼ��ؼ�漷��oc��Bfڼ�˼����ϵ��`����P   P   ��g���:"��~����t�;Kڼm�ȼ�g���Ȳ�,���_��ɰ���Ѿ��P��ڶ���ᵼ����m̼J�ݼP   P   u���'/��k8�l�7��-����MI����Ǽ�᭼�d��5ӓ�zҏ��d��V���mC��ڶ���˼$��ڽ
�P   P   O�F�p�U��|x������.n���K��H'�-��I�Լ�䬼���1)��������V���P��Bfڼ����*�P   P   9ȁ��R���J��݈ƽ�ƽ|ն�@P�����E������'M���̍��9~�����d��Ѿ����[�O>J�P   P   �\���JȽ�����,��3��v
���dŽY��._��� ��:輾쭼�̍�2)��zҏ���nc��$��@d�P   P   7����D��H�8���K��pK�]7�� ���(਽��m�P�$��:�'M�����5ӓ�ɰ����*)��*s�P   P   �Ų�:I ��^0�Epc��;��)��ȏ���Ga��.�H���H����m��� �����䬼�d���_���漬�$��s�P   P   N4���M �`T9��:~��'���0�����L��0r{�?�6�H��)਽._���J�Լ�᭼,����ؼz���d�P   P   �Q�����|0��b~�G ���Ҿ�����Ѿ����0r{��.���Y���E�-���Ǽ�Ȳ��xɼ�O�s�I�P   P   �Ɓ��vȽ?,�%�c��r���-Ӿ� ��E{����ѾL���Ga�� �dŽ���H'����g��"���I*��I*�P   P   �O�	��������H9�~���෾�J㾶 ��������ȏ��]7���AP����K�MI�m�ȼ�K����ʼ{]
�P   P   ���<q��ḽ���J�L�x؎�෾�-Ӿ�Ҿ�0��*���pK��v
�|ն�.n����<Kڼe��Jׯ���ܼP   P   ���/�������ǽ�+�J�L�~����r��H ���'���;����K��3��ƽ�����-��t����]&��e^��P   P   ����{�����9��n����ǽ����H9�&�c��b~��:~�Fpc�I�8��,�ވƽ}x��m�7����k���ӏ�A��P   P   ����h��������9������ḽ����@,�|0�aT9��^0�E�������J��U���k8�;"��)��������x�P   P   ��e������h��{����/��<q�	����vȽ����M �:I ����JȽ�R��G�p��'/�h�����������!e�P   P   �{ży̼�� %�-o�;�;�Z�b�����5&��G[���'���_��93��g���5�b�Y <�Fu�,���t�̼P   P   t�̼5T̼O7ռ��� ��di�|�+��1E��n^���r�M:~�iU~���r���^�ߞE���+����������ռP   P   ��8�޼�������`j���D��q�)���6�?@���C�{@�X7��$*���#���&�NF���P   P   ,����[�H��� �p�����������+J�i|���u������	��������&����P   P   Fu��H ���!����f��b�d]��^��M��� �I
 �,? �� ��� �� �ݥ�������#�����P   P   Y <�M0I�^EP�j�O���G�&Q:���)�8����u����k������9P��z����ݥ��	�����+�P   P   4�b���|�]v��t����熽F�z�``���B� �'�a��� �����n�ؼژԼ �ټ�z�� �����$*�ߞE�P   P   f����蛽,2��yz������#���a����<L[�4A4�6E�������ӼژԼ9P㼀� �u��X7���^�P   P   83��о���>ٽ�����ｫ�׽c������{o��*=��?�����n�ؼ��� ���{@���r�P   P   �_����ҽN�_���
"�4�!��� ��'нaᢽ<z�e@�����������,? �h|���C�iU~�P   P   �'��pE�����0���H�ϪQ�|�G��(/���!K޽���<z��*=�6E�� ���k�J
 �+J�?@�L:~�P   P   F[���O�g�Z}@���f�%r~���}���e�Z�>����!K޽aᢽ{o�4A4�a��u����� �����6���r�P   P   5&����ҽJ���@�k�r�!O��放�Ќ�,q�Z�>����'н���<L[� �'����M���q�)��n^�P   P   �����ٹ�	u���0�.Gg��r��f���e���Ќ���e��(/�� �c����󃽉�B�8���^����D���1E�P   P   Z�b���;�ٽ`Z��MI��1�KE��f���放��}�|�G����׽�a��``���)�e]������|�+�P   P   ;�;�N}�Ӟ��l�𽂱"��R��1��r��!O��&r~�ЪQ�4�!�ｌ#��F�z�'Q:��b�q�`j�di�P   P   -o�W�I��ꇽ�D��m����"��MI�/Gg�l�r���f���H��
"��������熽��G�f�� ��� ��P   P    %�C� ��	Q�2R���D��m��`Z���0��@�[}@��0�`����zz��u���k�O����I���漌��P   P   �����;i"��	Q��ꇽӞ��;�ٽ	u�J��g���N��>ٽ-2��]v��_EP���!�	[����O7ռP   P   y̼�߼���C� �W�I�O}����ٹ���ҽ�O�qE���ҽо���蛽��|�N0I��H ����9�޼5T̼P   P   ��2 ������"��7��	R�u	p��q��)�����W3��^����4��聇��(p�T*R�3�7�l�"�����P   P   ����˸�.���J"�B�1�]E�PQY��l��C|�Gr��yz���u|��	m�V�Y�/iE��r2���"�2�����P   P   ��^�����h�`d�r�"��4,�F�7�B C���M�8�T�C�W�((U�E�M�s�C��&8���,��U#�h��2��P   P   l�"��#���"�cY"�&�!��V"���#�F�&�u9+���/���3��36�jQ6�FC4��n0��,�	�'���$��U#���"�P   P   3�7�{�;�e�<�;�:���6�XD1��+��&��(#��2!��w ��� �v� �U� �z.!��+"�a$�	�'���,��r2�P   P   T*R�%9\�]�a�2Qa�!I[�I�P���C�e6�(x*��� �A��ѵ���g�N_�����+"��,��&8�/iE�P   P   �(p��聽Ω��a ��-A��($���%n���W���A���.�Q��Y�5M�|���N_�z.!��n0�s�C�V�Y�P   P   聇��ݗ�����HK������a:��c���}0��@bj��K��>2��l�x(�P+�|�g�U� �FC4�E�M��	m�P   P   �4���f��qUý?�ҽ~#ؽҽ½lޫ�_���>hy�ܕR�XJ4��H�x(�5M���v� �jQ6�((U��u|�P   P   ]����辽.9߽T���)���f�4���?�ݽ|����߀���T�XJ4��l�Y�ѵ��� ��36�C�W�yz��P   P   W3��p�Ƚ�@�˞�?7��z!�q��T���1��ƽyN���߀�ܕR��>2�Q��A���w ���3�7�T�Gr��P   P   ���Y�Ƚ����:W���-�n�:��:��-��O�c����ƽ�>hy��K���.��� ��2!���/���M��C|�P   P   )��,��a��e��r4��2J��1R���I�Y�3��O��1�|��_���@bj���A�(x*��(#�u9+�B C��l�P   P   �q���y��i߽����.�_\J�MA[��[���I��-�T��?�ݽmޫ�}0����W�e6��&�F�&�F�7�PQY�P   P   u	p�i�����ý�w��.��xa;���R�MA[��1R��:�r��4���½c����%n���C��+���#��4,�]E�P   P   �	R�����K���Pӽ)�R"�xa;�`\J��2J�o�:��z!��f�ҽa:��($��I�P�XD1��V"�r�"�B�1�P   P   �7�4j\�����y۬���ؽ)�.���.��r4���-�@7�*��#ؽ����-A��!I[���6�&�!�`d��J"�P   P   ��"�<�;�T(b�V���y۬��Pӽ�w������e�:W�̞�U���?�ҽHK��a ��2Qa�;�:�cY"��h�.��P   P   ��� ,#�,=�T(b������K����ýi߽�a������@�/9߽qUý����Ω��^�a�e�<���"���˸�P   P   2 �� ,#�<�;�4j\����i����y��,�Y�Ƚq�Ƚ�辽�f���ݗ��聽%9\�{�;��#�^����P   P   �u&�^�(�/0��l<��(M��a���x����5�����b���\
��+!�����-�x���a�uJM�%�<��I0���(�P   P   ��(���(�p,�^�2� @<���H�	�W�
�g��^v�>����:��\>�������v���g�X�LI���<���2��>,�P   P   �I0�XW/��0��p2�}a6���<��1D�TM��]V�VZ^���c�c�e�?d���^�e�V�L�M��D��$=�z�6���2�P   P   %�<�
x<��O<�� <���;�yP<���=��*@�aC���F�t�I� �K���K��JJ�`zG�6D��A���>��$=���<�P   P   uJM���O���P���O�ޑL�SVH�.�C�D�?�=�B);��v:�p7:�<V:�߄:�;��<���=��A��D�LI�P   P   ��a���i�2�m�B�m���h���`���V��DL��B���:��:5��v1�ޱ/��/���1�Y 6��<�6D�L�M�X�P   P   -�x�惽I�-���ࠈ��T���mw��7f�
/U���E���9�N$1�e�+�~�*�.p,���1�;�`zG�e�V���g�P   P   ����������#���q������_C��5����t���\�ڰH�SK9��$/�]N*�~�*��/�߄:��JJ���^���v�P   P   +!��4v��g���:=������Yɼ�l߱�ca��^����b�JJ��;9��$/�e�+�ޱ/�<V:���K�>d����P   P   \
��p�����Ž}W׽�2�
���ֽV�Ľ�d�����_����c�JJ�SK9�N$1��v1�p7:� �K�c�e�\>��P   P   b���4���b�ҽ��콣���ɉ�u!��V�뽠�ѽ�!���.��_���b�ڰH���9��:5��v:�t�I���c��:��P   P   ���&�����׽G���
����K��h�	��r���Aֽ�!����������\���E���:�B);���F�VZ^�>���P   P   5��������ҽ]���@���y�"�*�}T��r����ѽ�d��^��t�
/U��B�=�aC��]V��^v�P   P   ���v�����Ž��콃 
�G��U$�B�#�*�h�	�V��W�Ľda��5���7f��DL�D�?��*@�TM�
�g�P   P   ��x�R���鲽��׽�3��^��AA�U$�"�K��v!���ֽl߱�_C���mw���V�.�C���=��1D�	�W�P   P   �a���uŝ����b��x��^��G���y����ɉ�
��Zɼ������T����`�SVH�yP<���<���H�P   P   �(M�_�i�{"��M	�����c���3��� 
�A��
������2ὐ���q��ࠈ���h�ߑL���;�}a6� @<�P   P   �l<��P��'n���M	�������׽���^���G������~W׽:=��#���-���B�m���O�� <��p2�^�2�P   P   /0�(�<��JQ��'n�{"��uŝ��鲽��Ž��ҽ��׽c�ҽ��Žg�������I�2�m���P��O<��0�p,�P   P   ^�(��l/�(�<��P�_�i���R��v�������&���4���p���5v�����惽��i���O�x<�XW/���(�P   P   z>��@��ZF� P�C_]��Im�z�~����`���^������a��Np������~�Uym���]�<P��F��@�P   P   �@�̀@��C��UH��+P��8Z��e�s�q���|�Ă�I'���2���߂�N"}��r��.f�?�Z�ÈP�t�H�$GC�P   P   �F���E��TF��BH��K�?~P�9�V�[�]�w|d�Śj�ξn�|Lp���n���j���d�{^�Y&W�� Q�
*L�t�H�P   P   <P��9P��P���O���O��eP��ZQ�5cS���U��sX�ٷZ�_\��/\��[���X�daV��T�R�� Q�ÈP�P   P   ��]�8�_��Z`�pc_���\�'�Y�TKV�u/S�D�P��BO�g�N�):N�1kN�?{N���N���O�Y�Q��T�Y&W�?�Z�P   P   Uym��Is�(Cv��v�m�r�l�l��e�N]��TU�� O�%UJ��(G�t�E��E�+�G��K���O�daV�{^��.f�P   P   ��~�����>����ĉ��`��������}���p�|�c�9�W��N��F���B�V�A��7C�+�G���N���X���d��r�P   P   ���ِ�Γ���:��L���(���7���X���{�[ui���Y���M��bE�B\A�V�A��E�?{N��[���j�N"}�P   P   Np��bכ�~������)��,`���好*��������[m���Z��M��bE���B�t�E�1kN��/\���n��߂�P   P   �a��Qq���z���U��G�ŽʍŽ�˾�{���ہ���n��KP��[�n���Z���M��F��(G�):N�_\�|Lp��2��P   P   ���� ���l��z?ͽ�ؽ��ܽrؽ��̽2}���"�����KP��[m���Y��N�%UJ�g�N�ٷZ�ξn�I'��P   P   �^���%������4ս�����m� ���/Խਾ��"���n�����[ui�9�W�� O��BO��sX�Śj�Ă�P   P   `��Jr���q��ս$��~K��/������eH��/Խ2}��ہ������{�|�c��TU�D�P���U�w|d���|�P   P   ����՛�Ǒ���bͽgB��e����������� �彁�̽{���*���X����p�N]�u/S�5cS�[�]�s�q�P   P   z�~��֐�ٝ��\���� ٽt���������/����m�rؽ�˾��好�7����}��e�TKV��ZQ�9�V��e�P   P   �Im����O���Dﭽ�ƽ�Uݽt���e��~K������ܽʍŽ,`���(������l�l�'�Y��eP�?~P��8Z�P   P   C_]�jLs������x�������ƽ� ٽgB�$�����ؽG�Ž)��L���`��m�r���\���O��K��+P�P   P    P���_�({v����x��Dﭽ\����bͽս4սz?ͽ�U�������:���ĉ��v�pc_���O��BH��UH�P   P   �ZF�fDP�o�`�({v�����O���ڝ��Ǒ���q�������l���z��~��Γ��>���(Cv��Z`��P��TF��C�P   P   �@���E�fDP���_�jLs�����֐��՛�Jr���%��� ��Qq��bכ��ِ������Is�8�_��9P���E�̀@�P   P   l�Q��S��W�&Y_�_}i�ɡu�5\��������������鑽������������o��o�u��i���_���W��%S�P   P   �%S�]S�m.U�'_Y�^^_�g�I�o���x�æ���Ӄ�B���à���惽yŀ��@y�Z=p��cg���_���Y��OU�P   P   ��W��HW���W��PY�\�U�_���d�s�i��	o���s��v���w���v���s�jo�4:j��e�-I`��r\���Y�P   P   ��_�a_��K_�+:_��=_���_�^�`��
b���c���e�%|g��dh��{h���g�@f�?xd���b��9a�-I`���_�P   P   �i�:k���k�c�j��8i���f�1Hd�}�a�Z`���^��(^���]���]��^�.�^�fr_���`���b��e��cg�P   P   o�u�o0z�h_|��8|���y�//u��eo�K^i�ڜc���^���Z��gX�d5W�KW���X��T[�fr_�?xd�4:j�Z=p�P   P   �o��s������������y�����2Cx��cn��Te��]��>X���T���S��:U���X�.�^�@f�jo��@y�P   P   �������璽h����v��Ś���Y4��^0����r�o�f�(b]���V���S���S�KW��^���g���s�yŀ�P   P   �������>���ќ���E���\���"��Og��i���B����u�p�g��]���V���T�d5W���]��{h���v��惽P   P   �������쇦�"���.岽xò��6��@����h��-�C���Ҿv�p�g�(b]��>X��gX���]��dh���w�à��P   P   �鑽t`��7����߷�����4½�I���b��5�������5��C�����u�o�f��]���Z��(^�%|g��v�B���P   P   ���c��2������.ȽAν�ν��ǽSy���������-󏽃B����r��Te���^���^���e���s��Ӄ�P   P   ���������������P˽��ԽFKؽڳԽ��ʽSy��5����h��i��^0���cn�ڜc�Z`���c��	o�æ��P   P   �����񕽛���F���GȽ�
ս@ܽ��۽۳Խ��ǽ�b��@���Og��Y4��2Cx�K^i�}�a��
b�s�i���x�P   P   5\��R��y�������7����wν'sؽ@ܽGKؽ�ν�I���6���"�������eo�1Hd�^�`���d�I�o�P   P   ɡu��l������f����"���½�wν�
ս��ԽAν�4½xò��\��Ś��y��//u���f���_�U�_�g�P   P   _}i�}&z�{/������Z����"��7���GȽ�P˽.Ƚ���.岽�E���v��������y��8i��=_�\�^^_�P   P   &Y_�>7k�x|��7������f�������F����������߷�"���ќ��h�������8|�d�j�+:_��PY�'_Y�P   P   �W��]_�8�k�x|�{/������y�����������2���7���쇦�>����璽���h_|���k��K_���W�m.U�P   P   �S�^BW��]_�>7k�}&z��l��R�������c��t`�����������s��o0z�:k�a_��HW�]S�P   P   T`�4ia��e�K�j���r�Z�{����^���@��~ʍ������Ӎ��H��;u�� ӂ�/ |� �r��k��e��a�P   P   �a�xoa�c�Rf�4k�4�p���w��O~�i6��[���NɅ�M˅�����AU��L�~�[�w�.Kq��Ok�`�f�r-c�P   P   �e�p�d�� e�}@f��Lh�Qk���n�m�r�2�v�+z�x|��T}��|��_z��.w�PDs�rYo��k�v�h�`�f�P   P   �k��j��j���j���j�<8k��	l��m�9jn�9�o�k�p�/�q���q�):q��p�1�n���m���l��k��Ok�P   P    �r�x�s��Gt���s�5�r��p���n���l��pk��sj�
�i���i��i��i�LCj���j� l���m�rYo�.Kq�P   P   / |�X�~��Z���N��0�~��|{�9w�d�r�G(n��cj��mg��fe��~d�Y�d�j�e�E�g���j�1�n�PDs�[�w�P   P    ӂ��ȅ�0���S�����
����z����}��gv��mo�&�i�lMe���b��b���b�j�e�LCj��p��.w�L�~�P   P   ;u���������9@���'���L��e����	���恽�y�~p�	Oi�4>d�7�a��b�Y�d��i�):q��_z�AU��P   P   �H������h����x�������N��{���WB���ӊ�6��%�{��,q�pi�4>d���b��~d��i���q��|�����P   P   �Ӎ���>��9������f���%z���؜��|��X��EQ��>z|��,q�	Oi�lMe��fe���i�/�q��T}�M˅�P   P   ����WH���m��.���D����������֨��������v>��EQ��%�{�~p�&�i��mg�
�i�k�p�x|�NɅ�P   P   }ʍ�W@���⢽r���,
������᷽�ĳ�/;���h������X��6���y��mo��cj��sj�9�o�+z�[���P   P   �@�����u������: ���L�������(��'���/;������|���ӊ��恽�gv�G(n��pk�9jn�2�v�i6��P   P   ^��d���X@��U7�����qa�����������(���ĳ��֨��؜�WB���	����}�d�r���l��m�m�r��O~�P   P   ����������*Ѣ�?^��d��z�����������᷽���%z��{���e����z��9w���n��	l���n���w�P   P   Z�{�����R���񐚽Y好�.��d��qa���L����������f����N���L��
����|{��p�<8k�Qk�4�p�P   P   ��r���~�����[��,ț�Y好?^�����: ��,
���D����������'�����0�~�5�r���j��Lh�4k�P   P   K�j�`�s�xc��Yl���[��񐚽*Ѣ�V7������r���.��9����x��9@��S���N����s���j�}@f�Rf�P   P   �e���j��Tt�xc�����R�������X@���u���⢽�m��>��h�������0����Z���Gt��j�� e�c�P   P   4ia���d���j�`�s���~��������d�����W@��WH������������ȅ�X�~�x�s��j�p�d�yoa�P   P   �hk�8zl��/o�ɋs��oy�!��*�������ԉ�󳋽pY��/���䉽���=����'���y�G�s��Ho���l�P   P   ��l��l���m��1p���s��#x�n)}�M���9�������ꅽ;酽����M��g)���c}�fx���s�1`p�-�m�P   P   �Ho��n��0o�<1p���q�at�6�v���y���|�D�([��n���2j���:��|��z�w�>Yt�|+r�1`p�P   P   G�s���s��s��|s�a�s�2�s�_�t�ku�{gv�vw��=x���x���x�xex���w�=�v�:�u��t�>Yt���s�P   P   �y�qlz�A�z��Hz��Ky�T x���v��Qu�NFt�&hs�K�r�Y�r��r��r��7s���s�W�t�:�u�w�fx�P   P   �'���O���ぽgځ��2��f��.�|�q�y��7v�
Vs�%q�V�o���n���n���o���q���s�=�v��z��c}�P   P   =����م�zJ������h-��E����r�����7D|��,w���r��zo�o]m���l�ߌm���o��7s���w��|�g)��P   P   ����`��1挽�;��Y.��t���k#��3ǆ�����đ~���w�DXr�w�n�Y�l���l���n��r�wex��:��M��P   P   䉽w���9��?����������������.��8����������a@x��Or�w�n�o]m���n��r���x�2j�����P   P   /���Cx��7�������$���!����X���c���!��v[�������Q��a@x�DXr��zo�V�o�Y�r���x�n���;酽P   P   pY��N��E����ݞ�ab��L���KB�������>����|������������w���r�%q�K�r��=x�([���ꅽP   P   󳋽-�����C��fB��_����悔���a����R����v[������đ~��,w�
Vs�&hs�vw�D�����P   P   �ԉ��v��G���C����������d���׫��t��a����>���!��8�������7D|��7v�NFt�{gv���|��9��P   P   ����r�����;ꞽ�K��S���.䮽�Ϯ��׫���������c���.��3ǆ����q�y��Qu�ku���y�M��P   P   *����V��6�������w������y��.䮽�d���悔KB���X������k#���r��.�|���v�_�t�6�v�n)}�P   P   !���Ӆ��댽����y���x������S������_���L���!�������t���E���f��T x�2�s�at��#x�P   P   �oy�'I��LI��kK������y����w���K������gB��ab��$�������Y.��h-���2���Ky�a�s���q���s�P   P   ɋs��Sz��끽�ć�kK����������;ꞽC��C���ݞ�����?����;������gځ��Hz��|s�<1p��1p�P   P   �/o��s�2�z��끽LI���댽6�����G������E���7����9��1挽zJ���ぽA�z��s��0o���m�P   P   8zl���n��s��Sz�'I���Ӆ��V���r���v��-��N��Cx��w���`���م��O��qlz���s��n��l�P   P   �t���t���v�&=z�͋~�Z����\���ֆ��ˈ��#��<����'���܈�=↽�s��\с�ç~�`Oz�}�v���t�P   P   ��t��t�ˣu�ܒw�w?z�P�}�Y����x��I���K���1����U���&��莂�$���_�}��mz��w�Ϳu�P   P   }�v��v���v��w���x�r�z�Q�|��~��c��~S��*偽�#����b��$���r�~���|�K�z��y��w�P   P   `Oz�� z�yz�-z��7z�'�z���z��u{�r7|�K�|�A�}�C�}�!~���}�D.}�Cm|�O�{��8{�K�z��mz�P   P   ç~�5�;���k~��u}�||�l{�ޥz��y�7�y�cy�$Vy�N�y��y��Az��{�O�{���|�_�}�P   P   \с�p���������͕��D�������X�~�=|�u�y�#x��w��zv���v��>w��`x��Az�Cm|�r�~�$���P   P   �s����������PF���چ��҅��F��U���J����|��oy���v��}u���t���u��>w��y�D.}�$���莂�P   P   =↽iH��&�����닽�ފ����묆��能g&��VQ}��-y��Mv���t���t���v�N�y���}��b���&��P   P   �܈�?#��ӎ�R�������p��H����틽P������C�����}�ty��Mv��}u��zv�$Vy�!~���U��P   P   �'���I������������c���１�����䉽=��� ꁽ��}��-y���v��w�cy�C�}��#��1���P   P   <����p�������������욽����~������]8���T��=���C���VQ}��oy�#x�7�y�A�}�*偽�P   P   �#��yu��k��� P��,�e���׆��n���� ��z��]8���䉽���g&����|�u�y��y�K�|�~S���K��P   P   �ˈ�D�������O������K���2���L}������� ���������P����能�J��=|�ޥz�r7|��c��I��P   P   �ֆ����Gܮ��<ɜ�퓠�Ҫ��͡��L}��n����~��１��틽묆�U��X�~�l{��u{��~��x��P   P   �\��_?���Ԏ�E���)��c���N���Ҫ��2���׆�����c���H�������F������||���z�Q�|�Y���P   P   Z���J�'���@�������c���퓠�K���e����욽�񕽸p���ފ��҅�D����u}�'�z�r�z�P�}�P   P   ͋~����p[����-����)��<ɜ�����,�����������닽�چ�͕���k~��7z���x�w?z�P   P   &=z�$"�����R��[���@���E���ܮ���O�� P���������R����QF������-z��w�ܒw�P   P   ��v�z�?����p'����Ԏ�G����k��������ӎ�&����������;�yz���v�ˣu�P   P   ��t���v�z�$"����J�_?�����D��yu���p���I��?#��iH������p���5�� z��v��t�P   P   J�z�� {���|���s���&̈́��������� ��HV�����g�������ۄ�9���c"���$��|��{�P   P   �{���z�A�{��'}��$�π����l�����������������������;{���-��8〽@M��@}���{�P   P   �|�;M|���|��!}���}��K�3k���<��M�������;���7�����	���~��YS������v��%~��@}�P   P   �$�B�����5�C�������IQ��_������怽뀽р�@���3h��*��/��v�@M�P   P   c"���P��q��7B������ǀ��c���
��e�3�Z�~���~�xi~���~���~�,;�3��*������8〽P   P   9�������냽D僽�w���Ⴝ���v*���E��k�~�9�}�Ȳ|�9L|��O|�|�|��}�,;�3h��YS���-��P   P   �ۄ�' ������ ��������ⅽɹ���S���偽�v���~���|�|�{��>{�)�{�|�|���~�@���~��;{��P   P   �����_������FL��4A��䓉��=���t��G���i��d���Sa~��*|��*{��>{��O|���~�р�	������P   P   g��*h���X��y������F���w>���=���燽�\����������+A~��*|�|�{�9L|�xi~�뀽�������P   P   ���������?q����9x��j\��[g��-ۋ�؈��ԅ�`������Sa~���|�Ȳ|���~��怽�7�����P   P   HV��i͌�9
������%T���蔽�E��A����ᏽ����w(���ԅ�����d����~�9�}�Z�~���;������P   P   � ���͌�(v��l����8��Ax��\s�����\���I������؈��\��i���v��k�~�3�_�����������P   P   ���� ���
��hǓ��ז�̘�q����ָ��\����ᏽ-ۋ��燽G����偽�E��e�IQ��M������P   P   ����xd��`���G���Z;��yј��G��>F������A���[g���=���t���S��v*���
������<��l��P   P   &̈́��W��WY��fy���Y������$����G��q���\s���E��j\��w>���=��ɹ������c�����3k�����P   P   �����0���;���������������yј�̘�Ax���蔽9x��F���䓉��ⅽ�Ⴝ�ǀ�C��K�π�P   P   s�����������O����������Y��Z;���ז��8��%T�������4A�������w�����5���}��$�P   P   ��fI���烽����O��;���fy��G���hǓ�l�������?q��y���FL�� ���D僽7B�����!}��'}�P   P   ��|�>�et���烽����0���WY��`����
��(v��9
�������X����������냽q������|�A�{�P   P   � {�A|�>�fI�����������W��xd��� ���͌�i͌���*h���_��' �������P��B�;M|���z�P   P   �
���'_���=���|���Ճ��=��`��������,���n���0��q���򌆽BG��_僽؇���K���d��]��P   P   ]��~�����ŕ���X��z:��!9��!7������������������D���A���J��,I��Oe������#��P   P   �d��S���^���[���Xo��X큽�������w���D能�����탽����x)��£��������2������P   P   �K���G��SE���@���U���i��Ќ��ѵ��6݁�����5���G��`I��tC�����Q���@Ɂ�A������Oe��P   P   ؇��8���z�������e{��y3���恽�����e��Q<��m��]��V�����D0���R��[���@Ɂ����,I��P   P   _僽zN�� x���p��~C��EɃ�y2�������؁��<��+����j��aG��VM���x��pՀ��R��Q���£���J��P   P   BG��
��j���ﱆ����n����)���(�����c���s��	k��������4���x��D0�����x)���A��P   P   򌆽@�������������͓������j���[���$�����9A��d�����VM�����tC������D��P   P   q���F�����fs��t���`i��g���=)��k�����j΃��/�����9A�����aG��V��`I���탽���P   P   �0��4P���.��K���f4��!6��r�����'0������ⅽ,ჽ�/�����	k���j��]���G���������P   P   �n��j튽�-�����X/��N���T#���򎽚���Ɗ��T���ⅽj΃�$��s��+���m���5��D能���P   P   �,���䊽5����ԏ�\����d��b��3o��o���>v���Ɗ�������[���c����<��Q<�����w�������P   P   �����N��!-��g؏�����1f���ד��^���ᑽo������'0��k�������؁��e��6݁�������P   P   `����?��-��z	��A����h��tH��e=���^��3o�������=)���j���(����������ѵ������!7��P   P   �=��]���D���5����4���g��F���tH���ד�b��T#��r��g�������)��y2���恽Ќ��X큽!9��P   P   �Ճ�
�����v��?��̞���g���h��1f���d��N���!6��`i��͓��n���EɃ�y3���i��Xo��z:��P   P   �|��2H������J������?���4��A�������\���X/��f4��t���������~C��e{���U��[����X��P   P   �=�������s��~���J��v��5���z	��g؏��ԏ����K���fs�����ﱆ��p�������@���ŕ��P   P   '_���C��U����s���������D���-��!-��5����-���.���������j��� x��z���SE���^�����P   P   ��HT���C������2H��
��]����?���N���䊽j튽4P��F��@���
��zN��8����G��S��~��P   P   �Y��`���^끽՟��|r��e���l���Y��]�������̇����/$��Ha��>w���n��1���5�����������P   P   ����G���멁����Ɲ���K�����-���.S��4ƅ������� х�;Z��Ƅ�k��;V��y������x���P   P   �����災쁽���T�������������탽EC��'{�����@���8L��r���񓃽�*��[Ă�$a�����P   P   5���C���������������ȱ���͂�[����.���B���Z��{]��.K���;�������������[Ă�y���P   P   1�������}������cp���E������Ⴝ�����������om���r���u�����������ւ������*��;V��P   P   �n��U���iꄽ�䄽����]������~��9��-����9��M���*ց�oہ�����J���������񓃽k��P   P   >w��w�� o��a���ld��*��� c��Y���b����&���t������𩁽����*�����������;��r���Ƅ�P   P   Ha��aC�����N���O��{⇽�2��CG���>���2���:��Se���΁���������oہ��u��.K��8L��;Z��P   P   /$���X��=V��
)-���뉽�C���D�����t����c��BK��>_���΁�𩁽*ց��r��{]��@��� х�P   P   ���� ���q��0q��,����苽�c���a��0������n텽hx��BK��Se������M���om���Z��������P   P   �̇������%������d��L����Z���s�����Vx��T���n텽�c���:���t���9������B��'{�����P   P   ���������s��a���@���㎽ݎ��9�������b��Vx������t����2���&��-��������.��EC��4ƅ�P   P   ]������#���������r����叽p��������������0������>��b���9����������탽.S��P   P   �Y���R���t������/E��k����O�� J��p����9���s���a���D��CG��Y���~���Ⴝ[����-���P   P   �l��?��)R��Bm��Ce���뎽㏽�O���叽ݎ��Z���c���C���2�� c����������͂������P   P   e��^���Q���M����w����뎽k���r����㎽L����苽�뉽{⇽*���]���E��ȱ�������K��P   P   |r��&����i���P���7�����Ce��/E�������@���d��,���)-���O��ld������cp�������T��Ɲ��P   P   ՟�������넽/����P��M�Bm���������a�����0q��
�N��a����䄽������������P   P   ^끽{��������넽�i��Q���)R���t���#���s���%���q��=V���� o��iꄽ}�������쁽멁�P   P   `����䁽{�������&���^���?���R�������������� ���X��aC��w��U�������C����災G���P   P   x���ķ���	��9���x!���ꄽ	����F���҆��+��F��s/��CՆ�6K��_���c1�����c��?���P   P   ?���9����܂�3��X��������6��䒅�$ۅ����{����������d��o���S"������:������P   P   c������G��R5���Z������E탽�9��8��������焽J���"ꄽwǄ�t���oD������y���fh��:��P   P   ���q���腃�Ԋ������ݞ��Y�������Wڃ�3C��������*
�������僽�Ѓ�����y�������P   P   1���:��L���4���#��
��H샽���:���݁��%x���m���f��ir��:�����������Ѓ�����S"��P   P   cT���F���D�����脽΅��5��$փ��}��4=���������q�������I�������僽oD��o���P   P   _���t��rI���d��?D��@��}����������烽1v��I
��*˂�\���Gт����:�������t���d��P   P   6K�������n��V���]����b����;������������Le��U�پ��\���q���ir��+
��wǄ�����P   P   CՆ�Z���?j��t㈽�	���ڈ�}`�������Æ��υ��Մ������a��U�*˂������f�����"ꄽ����P   P   s/���S���<��b߉�e>���3���ى�b.���A��g��� ��g�������Le��I
������m�����J���{��P   P   F��y����ĉ�W����:��uq���:������:�������.��� ���Մ����1v��4=��%x��C���焽���P   P   �+������5㉽����틽�^�� [���拽����؉����g���υ����烽�}��݁��3����$ۅ�P   P   �҆��K���ŉ����)���ό����fȌ��"�����:����A���Æ���������$փ�:���Wڃ�8���䒅�P   P   �F�������8��6�����ӌ��P���T��fȌ��拽����b.�������;�����5����������9��6��P   P   	���k����i��<㉽=���a��9���P����� [���:���ى�}`���}���΅��H샽Y���E탽���P   P   �ꄽa���f���ވ�eA���o���a���ӌ��ό��^��uq���3���ڈ��b��@��脽
��ݞ��������P   P   x!��~��,H��!���;��eA��=���)���틽�:��e>���	��]���?D������#�������Z��X���P   P   9����4���D���g��!����ވ�<㉽6���������W���b߉�t㈽V����d���D���4��Ԋ��R5��3��P   P   �	��y����H���D��,H���f���i���8���ŉ�5㉽�ĉ��<��?j���n��rI���F��L��腃�G���܂�P   P   ķ��!���y����4��~��a��k��������K������y����S��Z�������t��T���:��q�������9���P   P   6��������܃�t1��ŵ��x2�������:��Ι���Ն�����nچ������D�����}9������}8��7݃�\���P   P   \���d���NÃ��䃽�<��닄�g��]��h����腽\�����!酽���X_��9���c���A��3KÃ�P   P   7݃�8փ�ۃ��烽����K��K{������넽���=��J>���?�� ��;􄽰Ą������R���$��3P   P   }8���?��$?��-4��v:��%F���X��mg���v��񈄽����ʘ��U���&���͎����s���c���R��A��P   P   ����$�������ַ��X���𐄽Pw��qk��FP���<��'��� ��s"���$���/��NG���\���s������c���P   P   }9���g��oo��o��,`���0���4����s���7�����Tჽu׃��׃��惽���NG����Ą�9���P   P   �������?���W���;������j���lV���ℽ:����*��|ჽ������� ����惽�/��͎��;�X_��P   P   �D����������8���2��Y���B���f7�����1��l���f��Y҃�?��������׃��$��&��� �����P   P   �����@��S������6,���������4��J����م� 6������[��Y҃����u׃�s"��U����?��!酽P   P   nچ�+����U���ۈ�������XՈ�FH�������̆�|���5������f��|ჽTჽ� ��ʘ��J>�����P   P   �����ᇽ�����b��dЉ�*�4Ή�^V��|���UՇ�V톽|��� 6��l����*�����'�������=��\��P   P   �Ն�7���	ڈ�G���eJ������+����?��d���?ʈ�UՇ��̆��م�1��:����7���<��񈄽���腽P   P   Ι��ԟ������C����q���� ��o��k��d���|�������J�������ℽ�s��FP���v��넽h���P   P   �:���?���N���_��EF�������D���G��o��?��^V��FH���4��f7��lV��4���qk��mg�������]��P   P   ����Ӧ������݈��Ӊ�b���k(���D�� ��+���4Ή�XՈ�����B���j����Pw���X��K{��g�P   P   x2��������F��������b��������񊽕���*������Y��������0��𐄽%F���K��닄�P   P   ŵ���c��;���;��X$�����Ӊ�EF���q��eJ��dЉ����6,���2���;��,`��X���v:������<��P   P   u1��D���jh���V���;��F��݈��_��C���G����b���ۈ����8���W��o��ַ��-4���烽�䃽P   P   �܃�D:��ǽ��jh��;�����������N������	ڈ������U��S��������?��oo������$?��ۃ�NÃ�P   P   ����i҃�D:��D����c����Ӧ���?��ԟ��7����ᇽ+����@����������g��$����?��8փ�d���P   P   �-��kD��
o������*
��g��hՅ�'#��r��领�F���٣��.x��E'���Յ��n�����@����l���G��P   P   �G��I��\��耄�����;����K�����������m ��w �������������ES�������Ä����X`��P   P   �l���d���j��い�B���c���섽���(7��CZ��Ei��Xq�� n��4]��f?�����p턽YǄ�~������P   P   @���Ы����������q���غ��V˄�Z΄�-ۄ��������k����񄽂愽�ք�Wф�YǄ��Ä�P   P   ���������6���������愽,˄�̻��ڴ��ʣ��u���*������a���Ը���Ą��ք�p턽����P   P   �n��g���+���Ȕ�������c��N��h���݄�䰄�����"s���^���a���v������Ը���愽���ES��P   P   �Յ�|��l/��`.���+�����(̅������2���섽6���Cr���P���C��CU���v��a�����f?�����P   P   E'�������ǆ�U熽�߆��ņ��y�����G����R���ꄽ����]��mB���C���a�����k���4]������P   P   .x��F솽�G��]w��
���~t��'<��ㆽ�o���녽�b����������]���P���^��*����� n������P   P   ٣��),���������S2��:6��s�������M#��J���(����e����������Cr��"s��u������Xq��w ��P   P   F����Y����m��4���i҈������k���臽uJ��m���(����b���ꄽ6�������ʣ���Ei��m ��P   P   领�&S�� ��ڢ������?���?���	��ڟ��6��uJ��J����녽�R���섽䰄�ڴ���CZ����P   P   r���/��Q뇽ͦ���,��_���x���Q���j"��ڟ���臽M#���o��G����2���݄�̻��-ۄ�(7������P   P   '#���ꆽ=���~n�����ʁ���ǉ���Q����	���k������ㆽ�������h��,˄�Z΄�������P   P   hՅ��|���@��� �����y?����ǉ�x����?������s���'<���y��(̅�N���愽V˄�섽�K��P   P   g��� ���ņ�b|��*3��hو�y?��ʁ��_����?��i҈�:6��~t���ņ�����c������غ��c���;���P   P   *
��ބ���*���ᆽs���*3���������,�����4���S2��
����߆��+��������q���B�������P   P   ����c��֘���+���ᆽb|��� ��~n��ͦ��ڢ���m�����]w��U熽`.��Ȕ��6������い�耄�P   P   
o������	��֘���*���ņ��@��=���Q뇽 ��������G���ǆ�l/��+�����������j��\��P   P   lD��Ic������c��ބ��� ���|���ꆽ�/��&S���Y��),��F솽����|��g������Ы���d��I��P   P   g�������ڄ���HA��*���oׅ����~E���m��jw���k���M��-���܅�����~C������܄����P   P   ���J���ʼ���愽���F���l������-ۅ��녽������%J؅�Ѧ���p���H�����섽�Ą�P   P   �܄��߄�R܄��焽�񄽛���2���H���u������J�������p���J���nw��cP���5��Z��S����섽P   P   ���	
��Y��
��h��)��b���(���2��'0���8���?���:���=���9���4���0���$��Z����P   P   ~C��}N��:W��JN���A��W@��@5�� %�����1��9
��q������-
��������"���0���5���H��P   P   ����۩����������4���9���<j��LE���/������턽ބ�Մ��ڄ����C����4��cP���p��P   P   �܅������K����F���օ�����t��1��L���܄�������������������9��nw��Ѧ��P   P   -���X��������������u~��TS������Ӆ�4{��+6��9���ф�7������ڄ�-
���=��J���J؅�P   P   �M��W���#膽q��{.��Z���ᆽ�����D��A酽����A6�������ф�����Մ������:��p���%P   P   �k���ކ�.7���s�����䛇�Uo��.6��MԆ�"b��� ��i���A6��9���܄�ބ�q���?���������P   P   jw�����j��=���Y������������b��/򆽤k��� ������+6��L���턽9
���8��J������P   P   �m������s��e函�6���f��:f���:��iڇ�[u��/�"b��A酽4{��1�����1��'0�������녽P   P   ~E��5܆��e������5K����������2����H��iڇ��b��MԆ��D���Ӆ��t���/������2���u��-ۅ�P   P   ��������;������):��	�������`���2����:�����.6������������LE�� %���(���H������P   P   oׅ�X���↽Ss��n����j��f�����������:f����Uo���ᆽTS���օ�<j��@5��b���2���l��P   P   *���������h��Ӛ��5���j��	��������f�����䛇�Z��u~��F��9���W@��)������F��P   P   HA���������t���T4��Ӛ��n���):��5K���6��Y������{.��������4����A��h������P   P   ���I��u������t���h��Ss����������e函=����s��q������K������JN��
���焽�愽P   P   �ڄ����KR��u�����������↽�;���e���s���j��.7��#膽����������:W��Y��R܄�ʼ��P   P   ����ۄ�����I��������X������5܆�����󆽣ކ�W����X�����۩��}N��	
���߄�J���P   P   v��,��!��3G��+{��@����؅����4��
J��U��M��V3��B��]܅�䩅��~��rI���#�����P   P   ���l��h���.��H���m��א��N���	ԅ��腽���������ꅽم�������	s���M���.�����P   P   �#��0���#���-���?��jW�� `��8���ԇ������n���v���߮��&���7��������i��WW�� F���.��P   P   rI��kO��~H��I���E���T��jM���T���^���_���r���g��k���p��ae��b��U[���R��WW���M��P   P   �~���{��Go���w�����Jm���d���X���L��]H��VC���7���;���<��xA���P���Q��U[���i��	s��P   P   䩅�����ͺ��»��	����������;~���[���I���6�����o������$���7���P��b���������P   P   ]܅�A�������!��C����Vڅ�ڹ������]���@��M��8�����c���$��xA��ae��7������P   P   B���;��]X��n���o���S���7��r���х����o���8��P������������<���p��&���م�P   P   V3��`n��F�������`���������Ok���-���䅽����1c���8��P��8��o���;��k��߮���ꅽP   P   M��嗆��Ԇ���	�����#��φ�u���:J����/���1c���8��M������7���g��v�������P   P   U��
���{���s8���a���k��#a��5���������ZM���򅽶���o���@���6��VC���r��n�������P   P   
J�������	��:W�����^�������)����T��^�����:J���䅽���]���I��]H���_�������腽P   P   �4��咆�O����T������Ǉ��Շ��ć�Ǜ���T������u����-���х������[���L���^��ԇ��	ԅ�P   P   ��m��ц��5�������ȇ�H퇽`��ć�)���5��φ�Ok��r��ڹ��;~���X���T��8���N���P   P   �؅�~;��R������Eb��o���*ԇ�H퇽�Շ�����#a��#�������7��Vڅ������d��jM�� `��א��P   P   @�����4U�����>���j��o����ȇ��Ǉ�^����k����������S�������Jm���T��jW���m��P   P   +{��B�����tp����>��Eb�������������a��	��`��o��C��	�������E���?��H��P   P   3G���~������� ��tp���������5���T��:W��s8��������n���!��»���w��I���-���.��P   P   !���G��:q��������4U��R���ц�O����	��{����Ԇ�F���]X�����ͺ��Go��~H���#��h��P   P   ,������G���~��B�����~;��m��咆�����
���嗆�`n���;��A��������{��kO��0��l��P   P   U9���F���U��nm��ʐ�������߅������ �� -���1��+2��N������݅��������r��QS���L��P   P   �L��F���U��B\��do��ڄ��%���&Å��х��������؅�T���������|o���]���V��P   P   QS���O��0V��Z��}j��_y�����r���ã�������������뺅�ٹ������B��������u��pr���]��P   P   r��Yr��[q��dn��mp��s���y������V���'������������������֑�� ������W���u��|o��P   P   ����F���ʤ��k���O����������������t��s��Ah���g���w���g��wl��}u��v�������������P   P   ��� �Kǅ��ʅ�����R�������皅����(v��jd���]���U��8N���a��eh��}u�� ���B�������P   P   ݅�6���������������6ۅ���������#���vh��+^���W���H��\���a��wl��֑������T�P   P   �����#���?���B���>���>��Q������ԅ�ɷ������ob��]S��CB���H��8N���g������ٹ���؅�P   P   N��tJ��$i����������,���Ai��ME������酽����Ҕ���v��]S���W���U���w�����뺅��P   P   +2��g������[����ˆ�n̆���������a���.���굅�Ҕ��ob��+^���]���g������������P   P   �1���p�����P�������k��"���qކ�����g���1�����������vh��jd��Ah������������P   P    -���l�������򆽵��95��4�����􆽊����g���.���酽ɷ��#���(v��s��'�������P   P   � ��e���������&��,J��mT��hL��^ ��������a�����ԅ���������t��V���ģ���х�P   P   ����<G�������ކ�r��N��*_���c��hL����qކ����ME����������皅���������r���&Å�P   P   �߅�@���m��f��������0��]X��*_��mT��4��"�������Ai��Q��6ۅ����������y�����%���P   P   ����F�K?��.��'Ά�����0��N��,J��95��l��n̆�,����>����R�������s��_y��ڄ��P   P   ʐ��~������SC�����'Ά�����r���&����������ˆ������>���������O���mp��}j��do��P   P   nm��ݛ��ʅ�P ��SC��.��f����ކ������P���[��������B�������ʅ�k���dn��Z��B\��P   P   �U��0n������ʅ����K?���m��������������������$i���?�����Kǅ�ʤ��[q��0V���U��P   P   �F��zT��0n��ݛ��~���F�@��<G��e���l���p��g��tJ���#��6��� �F���Yr���O��F��P   P   Wg���m���|��E���\��������ۅ�E􅽐�������� ��v�������ޅ�2ą��������U���dm��P   P   dm���t���i������Ǘ�����������ʅ� ᅽ�߅������텽�兽�ⅽ�Ʌ�����D���R���ʃ���k��P   P   U�������I���	�����������G���隅�N�������9���l˅�!�������
���
���}���斅�$���ʃ��P   P   ����=���膅����/��������������ə��ݝ������Û��՚�����������s���B���斅�R���P   P   ����������U��� ���ɥ��5���t���Ȗ�������������ք����������������s���}���D���P   P   2ą��ƅ��Յ��Ѕ��ǅ� �����-�������/���q}���y���r���r���y������������
�������P   P   �ޅ�셽A���������a�؅��ą�W������i����~��Kg��~s���l���y����������
����Ʌ�P   P   �������7���'��7)��E��.������Gޅ�j������Z���js��'p��~s���r������������ⅽP   P   v���-���?��(R���c��3T��@��[,�����������������|��js��Kg���r��ք��՚��!����兽P   P    ��<���`���u��愆�����r���`���8��#��2텽�ǅ�����Z����~���y������Û��l˅��텽P   P   ���^N��Ys��0�������P������!����t���K�����2텽������i���q}����������9�������P   P   ���L���w���������ˆ� ̆�����Ε���u���K��#������j������/������ݝ�������߅�P   P   ���?���p��{�������Dކ��↽�݆�"ņ�Ε���t���8�����Gޅ�W�������Ȗ��ə��N��� ᅽP   P   E�&*��wc��F������܆�O醽J䆽�݆�����!����`��[,�������ą�-���t�������隅��ʅ�P   P   �ۅ�'��@���q��䢆�̆�6熽O醽�↽ ̆����r��@��.���؅�����5�������G�������P   P   ����0l��5S��ȁ��q���̆�܆�Dކ��ˆ�P�������3T��E��a �ɥ�������������P   P   \����Ņ�����.&���e��ȁ��䢆��������������愆��c��7)���􅽏ǅ� ���/�������Ǘ��P   P   E��������ԅ�^���.&��5S���q��F���{�������0����u��(R���'�������Ѕ�U������	�������P   P   �|��툅� ����ԅ�����l��@��wc���p���w��Ys���`���?��7��A����Յ�����膅�I����i��P   P   �m������툅������Ņ�0'��&*��?��L��^N��<���-�����셽�ƅ����=��������t��P   P   ������������ŝ�����������م�$����1�����������>酽�څ�}Å�j���~����������P   P   ���� ���ď��.���>���n���e����˅��ԅ�8ᅽ�݅�߅�:ᅽ_ԅ��Ѕ������������ݕ�����P   P   �������e���j���ʗ������`���L���ٺ�����΅�`ʅ��х�8�N���*���گ��ʣ�����ݕ��P   P   ~���ä��Q����������f���Ɵ��Š��«��7�����������z�������	��������������ʣ�����P   P   j���,���ڳ��׹��|�������6�����������?�������f���f�������w���⣅��������گ������P   P   }Å��Ѕ��ͅ�Lȅ��х�Ką�����e�������Ԡ��*���䑅�#���W�����������⣅�����*�������P   P   �څ�V慽D酽\i녽W䅽�م��̅�ؼ������曅�􎅽̈��ϋ��򆅽����w���	���N����Ѕ�P   P   >酽����`	�������G�������셽N҅�ڼ������(���g���ޒ��ϋ��W�����������8�_ԅ�P   P   ����J���)��,/���%��c+���&��9�������ⅽn̅�x�������g���̈��#���f���z����х�:ᅽP   P   �����4���P���Q��:P���Q���2��������/߅��ą�x���(���􎅽䑅�f�������`ʅ�߅�P   P   ���%��+B��F^��iu���x��]v���^��-?��E(��Z���/߅�n̅�����曅�*������������΅��݅�P   P   1���(���K���n������:������������m��iG��E(������ⅽڼ������Ԡ��?���7�����8ᅽP   P   ��������?�� o��ϋ��f���5������������m��-?���������N҅�ؼ����������«��ٺ���ԅ�P   P   $t���4��/_�����`���Ы��Q������������^���2��9���셽�̅�e�������Š��L����˅�P   P   �م�� ��%��|Q���s������w���Ы��5�������]v���Q���&�������م�����6���Ɵ��`���e���P   P   �����ᅽ:��q.��vP���x������`���f���:����x��:P��c+��G��W䅽Ką�����f�������n���P   P   �����Ѕ�G텽5��H*��vP���s�����ϋ������iu���Q���%�����i녽�х�|������ʗ��>���P   P   ŝ��:���Uʅ��셽5��q.��|Q��/_�� o���n��F^���P��,/����\Lȅ�׹������j���.���P   P   ����8������Uʅ�G텽:��%���4���?���K��+B��4���)��`	��D酽�ͅ�ڳ��Q���e���ď��P   P   ����Ȇ��8���:����Ѕ��ᅽ� ��t������(���%����J������V慽�Ѕ�,���ä������ ���P   P   X���W���������������Ņ��ԅ��ۅ��셽��<��������텽�ᅽ�ׅ��Ņ����o���a���v���P   P   v���ᗅ�I���x�����������������ͅ�bۅ��څ��ޅ�Յ�΅�~ǅ�{���X����������l���P   P   a�������=����������ճ������컅�!����Ņ�
���2���]����Ņ�>���3������*���ɳ�����P   P   o���������������f���<���0���������������3���۹�����>���k�����������g���*�������P   P   ���1���清�����)����������޴��u���|���韅�F�����������$������������������X���P   P   �Ņ��ʅ�0˅�%ͅ��ą��Ņ�����ô��s���~�������إ��9���p�������������������3���{���P   P   �ׅ�=ޅ�O܅�
慽�߅�vׅ�)ԅ��Ņ�ܼ���������E���������[�������$���k���>���~ǅ�P   P   �ᅽ�酽y�������-���f���8݅�Eυ�+Å�����Þ��2���c������p�������>����Ņ�΅�P   P   �텽�������S�����=��������腽�Յ�6���2���1���2������9����������]���Յ�P   P   ����F	�������t.��1��- �����=�����ۅ�;���2���Þ��E���إ��F���۹��2����ޅ�P   P   <���^���)��w1��:���A��`5��|.��'����<��ۅ�6��������������韅�3���
����څ�P   P   ��5��o%��
3��'D��DO���P���@���8��K"�������Յ�+Å�����~���|��������Ņ�bۅ�P   P   �셽����*��E5���K���V���]��E\��4E���8��'��=��腽Eυ�ܼ��s���u�������!���ͅ�P   P   �ۅ��������r.���C��\��eX��s]��E\���@��|.��������݅��Ņ�ô��޴������컅���P   P   �ԅ��텽��#��6��|O��)a��eX���]���P��`5��- �����8)ԅ���������0�����������P   P   �Ņ��م�����`��E0��A��|O��\���V��DO���A��1��=��f���vׅ��Ņ����<���ճ������P   P   ����Bʅ��߅�t������E0��6���C���K��'D��:��t.�����-����߅��ą�)���f����������P   P   �������Lƅ��慽t���`��#��r.��E5��
3��w1�����S������
慽%ͅ�������������x���P   P   ����$���ܸ��Lƅ��߅�����������*��o%���)�������y���O܅�0˅�清�����=���I���P   P   W���ޞ��$�������Bʅ��م��텽�������5��^��F	�������酽=ޅ��ʅ�1�����������ᗅ�P   P   ܞ��y���D�������仅��ƅ��υ�/܅��ޅ��م�z兽l܅�ޅ��݅�҅��ȅ�W������������P   P   �������%���+���﵅�ظ��C����΅�@ׅ��Ѕ��ޅ�݅��Ӆ��օ�̅�ZÅ�:���������8���P   P   �������2���ᦅ�������������𵅽��������0����ʅ�6���Ną���������	���8���O������P   P   ����������B���ٷ��Ψ��ڲ��Y���c���Ӿ������׼�� ���#������������������8������P   P   W���4���j���ʵ��G���𺅽����9�������Ѯ��ڴ��|�����������󵅽	�����������	���:���P   P   �ȅ�DŅ��̅��Ӆ��ą��ą��ą�ٶ��-����������� �������H���K���7���	����������ZÅ�P   P   ҅�"ԅ��܅��؅�sم�9؅�D΅��ʅ�¾��[���.������a���ʯ��%���K���󵅽��������̅�P   P   �݅�߅� 腽煽����ꅽ�߅��م�)ׅ��Å�h������楅�����ʯ��H�������#���Ną��օ�P   P   ޅ�����r���������������	󅽱ᅽ�̅�������r���楅�a����������� ���6����Ӆ�P   P   l܅�b셽���p	�����.���	������څ�5م�c̅����������� ���|���׼���ʅ�݅�P   P   z兽�������	�� �����J��������R���Eꅽ5م���h���.�������ڴ������0����ޅ�P   P   �م�����s��p��:/��k,��~0��-�����(��R���څ��̅��Å�[�������Ѯ��Ӿ�������Ѕ�P   P   �ޅ����!��-���6��U5���7��1)���������ᅽ)ׅ�¾��-�������c�������@ׅ�P   P   /܅��>�����b-���3��z=���4���7��-����������م��ʅ�ٶ��9���Y���𵅽�΅�P   P   �υ��߅��􅽦��?!���*��C:��z=��U5��~0��J���	��	󅽧߅�D΅��ą�����ڲ������C���P   P   �ƅ��օ��酽q����������*���3���6��k,�����.������ꅽ9؅��ą�𺅽Ψ������ظ��P   P   仅���kօ�N䅽�������?!��b-��-��:/�� �������������sم��ą�G���ٷ������﵅�P   P   ���������Ѕ��ۅ�N䅽q���������!��p��	��p	������煽�؅��Ӆ�ʵ��B���ᦅ�+���P   P   D�������s����Ѕ�kօ��酽��>����s��������r��� 腽�܅��̅�j�������2���%���P   P   y������������������օ��߅�����������b셽����߅�"ԅ�DŅ�4��������������P   P   �����������䳅�z���i��������ƅ��Ѕ��݅�х�Tۅ��ԅ�Fą���"������Ͳ��k�������P   P   ����.���v�����������#���8���9��� �M̅�iŅ������υ���������޽��%���7���Ƴ��9���P   P   k�������ǫ���������+�������p���U���7����ȅ�G���%ȅ�������������(�������a���Ƴ��P   P   Ͳ�����洅�������������˶������2���-�������������B�������X�������޵������7���P   P   �������D�������������޹��^���᷅� ������������������c���ô��0�������(���%���P   P   "���ą�:��������ą��������1���^���;���+�����������������������ô��X�������޽��P   P   ��fʅ�(Ӆ�wʅ�{̅�2΅�QÅ�Y�������n�������:���Σ�����򧅽����c���������������P   P   Fą�+Յ�م�����j䅽م�Qх��ǅ�F�������n�����������Z��������������B�����������P   P   �ԅ��ޅ�C慽�䅽/녽�酽ㅽ�݅��Յ�rͅ��Ņ�����g�������Σ��������������%ȅ��υ�P   P   Tۅ�m煽rㅽE���
����񅽶��煽�����څ���������������:��������������G�������P   P   х�텽�煽n�_ ���������􅽌慽ꅽ�ԅ����Ņ�n�������+����������ȅ�iŅ�P   P   �݅�F텽
#������r��������s�����ꅽ�څ�rͅ�����n���;��� ���-���7���M̅�P   P   �Ѕ��兽mㅽ  �����������Z����s����慽�����Յ�F�������^���᷅�2���U��� �P   P   �ƅ��݅��煽 ���)��J������|��Z���������煽�݅��ǅ�Y���1���^�������p���9���P   P   �����х��䅽O�� ��"	���	���������������ㅽQх�QÅ�����޹��˶������8���P   P   i����υ�cم�l酽��:��"	��J������r������񅽣酽م�2΅������������+���#���P   P   z�������΅�G߅������� ��)���������_ ��
���/녽j䅽{̅��ą�����������������P   P   䳅�p���l����ʅ�G߅�l酽O� ���  ��#��n�E����䅽����wʅ��������������������P   P   ���J���v���l���΅�cم��䅽�煽mㅽ
�煽rㅽC慽م�(Ӆ�:���D�洅�ǫ��v���P   P   ��������J���p��������υ��х��݅��兽F텽텽m煽�ޅ�+Յ�fʅ�ą������������.���P   P   ]�������Y���Y������������ǅ��υ��ǅ��х��҅�SЅ�Ʌ�Jυ�
ʅ�����R���e���䬅����P   P   �������Ǭ��`��������������Կ���ȿ������"Ņ����'ą�����)�������ܴ����������P   P   䬅�<���Ū����������Ű�����"���׼��p���-���m���r���P���Ž��|�����������ﰅ�����P   P   e�������Ѳ���������;�������,���ѵ��ڳ��񷅽�������䴅�e���t�������E�������ܴ��P   P   R���.�����������5���A���K���"�������8���'���⭅�����⫅���������e���������������P   P   ����ݾ��&�������������������ڳ������ۭ������Ǳ��a�������0���ܴ������t���|���)���P   P   
ʅ��Å��Å��ͅ��ȅ������ȅ����Ƚ��W���(�������H���L�������0�������e���Ž������P   P   Jυ�,҅�E̅�#̅��Ѕ�%ǅ�Ѕ�υ�����¾��w���K���毅�׬��L�������⫅�䴅�P���'ą�P   P   Ʌ�ͅ�jх��م��ׅ��ׅ�ׅ��ͅ�dą��Å�����j�������毅�H���a�����������r������P   P   SЅ�Iׅ�ޅ��ᅽ�ᅽ3߅�)߅�&ޅ��Յ��Ѕ��Ņ�����j���K�������Ǳ��⭅����m���"Ņ�P   P   �҅�̅��兽#䅽텽+酽S腽c腽;υ��˅��Ņ�����w���(�������'���񷅽-�������P   P   �х�Jх��ۅ�|셽�����?셽�ꅽ�ۅ�;υ��Ѕ��Å�¾��W���ܭ��8���ڳ��p���ȿ��P   P   �ǅ��҅��煽�텽����?���l ��-����ꅽc腽�Յ�dą�����Ƚ����������ѵ��׼���P   P   �υ�υ��ޅ��腽Z녽�����������l ��?셽S腽&ޅ��ͅ�υ����ڳ��"���,���"���Կ��P   P   �ǅ� х�hӅ�a䅽�ⅽ���'�������?�����+酽)߅�ׅ�Ѕ��ȅ�����K��������������P   P   ����Å�ȅ�;Յ��䅽�腽�����������텽3߅��ׅ�%ǅ���������A���;���Ű������P   P   ����o����ȅ��υ� Յ��䅽�ⅽZ녽��셽䅽�ᅽ�ׅ��Ѕ��ȅ�����5�������������P   P   Y���y���ѹ��̅��υ�;Յ�a䅽�腽�텽|#�ᅽ�م�#̅��ͅ�����������������`���P   P   Y���Ǳ������ѹ���ȅ�ȅ�hӅ��ޅ��煽�ۅ��兽ޅ�jх�E̅��Å�&�������Ѳ��Ū��Ǭ��P   P   �������Ǳ��y���o���Å� х�υ��҅�Jх�̅�Iׅ�ͅ�,҅��Å�ݾ��.�������<�������P   P   .���\���䭅�'���笅�.���񶅽p����Å�f����ǅ�޾�������������������������ٯ��ꭅ�P   P   ꭅ�ʬ�����򫅽$���ذ������]���C���{�������0Å�+���������7�����������e�������P   P   ٯ��⭅� ���0���e���������������ᯅ�ð����Ӱ��b���ó��`���˱�����%�������e���P   P   ��������'�������-���&���P���[��� ������H�������%���²��ߴ��ӯ����������%�������P   P   �����������X���گ��k���ʰ��˺�����R�������(���򫅽l����������б�������������P   P   �������	���#������簅�Z�������쮅�%�������q���f���W������x������ӯ��˱��7���P   P   ����ṅ����i�����අ�������������ұ������S���������������������ߴ��`������P   P   ��������Ʌ����������Ņ�ֽ��T�����������2������'����������W���l���²��ó�����P   P   ����Å�ȅ�_х�[΅�,υ��ʅ�(�������J����������R���'�������f���򫅽%���b���+���P   P   ޾���Å�L̅�˅�IӅ��Յ�]̅��ą��ƅ��������Ĵ��������S���q���(�������Ӱ��0Å�P   P   �ǅ�ȅ��΅��Ѕ��օ��Ӆ��م�҅��Ѕ�?Ʌ�Wą���������1���������������H���������P   P   f����Ņ��Յ�ʅ�M܅��ۅ�؅��ۅ��΅�|ͅ�?Ʌ����J�������ұ��%���R������ð��{���P   P   �Å������Ӆ��̅�х�ׅ��Յ�օ�Ѕ��΅��Ѕ��ƅ�������������쮅���� ���ᯅ�C���P   P   p��������ǅ��υ�(ۅ�!݅��߅��兽օ��ۅ�҅��ą�(���T�����������˺��[�������]���P   P   񶅽?��� ȅ��̅�;څ��Ӆ��Յ��߅��Յ�؅��م�]̅��ʅ�ֽ������Z���ʰ��P�����������P   P   .���ճ���ȅ�΅�3օ��ׅ��Ӆ�!݅�ׅ��ۅ��Ӆ��Յ�,υ��Ņ�අ�簅�k���&�������ذ��P   P   笅�����ҽ�����ƅ�3օ�;څ�(ۅ�х�M܅��օ�IӅ�[΅����������گ��-���e���$���P   P   '���u���񼅽�����΅��̅��υ��̅�ʅ��Ѕ�˅�_х�����i���#���X�������0���򫅽P   P   䭅����ﮅ�񼅽ҽ���ȅ� ȅ��ǅ��Ӆ��Յ��΅�L̅�ȅ��Ʌ����	������'��� ������P   P   \����������u�������ճ��?������������Ņ�ȅ��Å�Å�����ṅ������������⭅�ʬ��P   P   ¥��ġ���������n���ٵ��^�������������0���������ش��y��������������������P   P   ������򨅽c���r�����������ɲ��γ�����������������u���䴅�G���a�������y���0���P   P   ���R���j���8�������2������m���D���ڭ��	������������������Χ��
���֨��y���P   P   ����>���󩅽妅�I���v��������������`���Y�������+�����������3���ʝ��L���
�������P   P   ���r��� ���3���Χ������㧅�<�������������¬���������������������ʝ��Χ��a���P   P   ����޵������Y��������������௅����������������{����������R�������3������G���P   P   y������̵��~���Ű��Ժ��f�������1�������5�������u���񥅽������������������䴅�P   P   ش��ӷ��z�������������������ѱ��U�������o�������y���e���񥅽�������������u���P   P   ���IÅ����� ����������������������]���n���%�������y���u���{������+�����������P   P   ���m�������	Å������Y�Å����W���;���E���%���������������¬�������������P   P   0���+ƅ�����B����˅��ą��Ņ��Å�
���!�����;���n���o���5����������Y���	�������P   P   �������eƅ��ͅ�҅��ͅ��Ѕ�rυ��̅��ƅ�!�W���]������������������`���ڭ�����P   P   ���+Å�&����Ʌ�Rօ�.ǅ�ԅ�"̅��Ӆ��̅�
���������U���1��������������D���γ��P   P   ��������ą�iÅ�҅�&Ʌ�[؅��Յ�"̅�rυ��Å�Å�����ѱ������௅�<�������m���ɲ��P   P   ^���D���=���v����˅�J΅�IՅ�[؅�ԅ��Ѕ��Ņ�Y���������f�������㧅�����������P   P   ٵ��ƹ��������]���Uȅ�J΅�&Ʌ�.ǅ��ͅ��ą������������Ժ����������v���2�������P   P   n���贅�E�������9�]����˅�҅�Rօ�҅��˅�����������Ű�����Χ��I�������r���P   P   ��������ů��,����������v���iÅ��Ʌ��ͅ�B���	Å� �������~���Y���3���妅�8���c���P   P   �������c���ů��E������=����ą�&���eƅ�������������z���̵������ ���󩅽j���򨅽P   P   ġ��|�����������贅�ƹ��D�������+Å����+ƅ�m���IÅ�ӷ�����޵��r���>���R������P   P   _���<���}�������]���F���ѥ�����������������?���*���ԫ���������ͪ��͢���������P   P   ���G���֣�����t���G���>���U���Q������P�����������𢅽쨅�ޝ��3���
���k������P   P   ����,���𧅽����ˠ����������١��m���W����������������/�����������*������k���P   P   ͢������	���נ�������񫅽���A�����������r������E���7���+���ƭ������*���
���P   P   ͪ������N���/���%���Ц������������)���s���(���塅�����墅����ѣ��ƭ������3���P   P   ����䦅�����$�������Т��^�������������I�����������?�������ר�����+�������ޝ��P   P   ���P�������"�����󥅽7���-���F����������������壅�!�������墅�7���/���쨅�P   P   ԫ��믅���������Y���I���M���N���>���E���c���͞����������壅�?�������E������𢅽P   P   *�������>�����������̯��>���[�������R���{���5���r���������������塅�����������P   P   ?���Y���[���������������I���v������İ������5���5���͞���������(���r����������P   P   �������"���(���N�����������}������򭅽�������{���c�����I���s�����������P���P   P   ��������Ѫ��Ҹ��z�������Q���ɮ��C�������򭅽İ��R���E����������)�������W������P   P   ����>�����������G����������J������C�������������>���F����������A���m���Q���P   P   ������������_�������n���r�������J���ɮ��}���v���[���N���-������������١��U���P   P   ѥ�����٭��P���
����������r�������Q�������I���>���M���7���^�������񫅽����>���P   P   F���٥���������������������n������������������̯��I���󥅽Т��Ц����������G���P   P   ]��������������N�������
�������G���z���N�����������Y���������%����ˠ��t���P   P   ��������1�������������P���_�������Ѹ��(���������������"���$���/���נ���������P   P   }����������1�����������٭����������Ѫ��"���[���>���������������N���	���𧅽֣��P   P   <���h��������������٥���������>�����������Y�������믅�P���䦅���������,���G���P   P   ~����������H�������d���N���礪����|���a���u�����������������������������\���P   P   \���#���얅�L���_�������������ɥ������M���ӥ��墅�Ҧ������T���u���T�����������P   P   ����ʗ����������Q��������������y���G����롅�
���>����������%������x�������P   P   ����͟��Ȝ������񜅽ԗ��M���@�������_���.����������ʟ��(���֖�������������T���P   P   ���Q���c���9�������/�������2���Ț�������������i�������"���Ԝ����������%���u���P   P   ����ף������D���L����������H���M���}���8���&���b���M���g�������Ԝ��֖������T���P   P   ������{���!���������M���A���@���J����������ϝ��v���t���g���"���(����������P   P   �������\���l�������t�������B���f���t���Y������՛��դ��v���M�������ʟ��>���Ҧ��P   P   ��������s���߮��礪�1���K�����������������D���	���՛��ϝ��b���i������
���墅�P   P   u���v�������̡�����%���~������0���󩅽������D����������&����������롅�ӥ��P   P   a������Ȳ�������������H����������<���D����������Y������8�������.����M���P   P   |�������U�������B���G���ૅ�ڴ��_�������<���󩅽���t���J���}�������_���G�������P   P   ���*�������ı����������8���U���e���_�������0�������f���@���M���Ț������y���ɥ��P   P   礪�Z���m�������鴅�����[�������U���ڴ������������B���A���H���2���@����������P   P   N���V���g���Ȥ��8������鉶�[���8���ૅ�H���~���K�������M����������M�����������P   P   d�������3���,���٩��q��������������G�������%���1���t����������/���ԗ��������P   P   ����Y�������	���٩��8���鴅�����B���������礪��������L�������񜅽Q���_���P   P   H���̠������"����,���Ȥ������ı����������̡��߮��l���!���D���9�����������L���P   P   ����h��������������3���g���m�������U���Ȳ������s���\���{�������c���Ȝ������얅�P   P   �������h���̠��Y�������V���Z���*����������v�������������ף��Q���͟��ʗ��#���P   P   d���ȕ��]�������-���И��ᙅ�&���B���S���}���ĕ���������악��������ɝ��`�������P   P   ��������ם�����`���3���$���e�������𘅽�������'���]���`����������D���C�������P   P   `�������o�������{���!��������������ٖ��#�������g���+�������曅�
����<���C���P   P   ɝ������隅�ћ������E�������:�����������������������Q�����������˕��9����D���P   P   ����������������/���$�������ܘ��1��������������Ő�����������������˕��
������P   P   ���%�������Y������虅�E���Ȗ�������������%���ؘ�����2���������������曅�����P   P   악��������y���������������֔������,������������������p���2��������������`���P   P   ����l����������������򑅽����&�����������ߗ��\���l��������������Q���+���]���P   P   ���������������$��������������\���n�������������\�������ؘ��Ő������g���'���P   P   ĕ������ԡ�����E���-���b�������М��딅�䛅�ښ�����ߗ������%������������������P   P   }���֠�����Y���e���"���ߣ���������u���p���䛅�����������������������#�������P   P   S���ݜ��񠅽񜅽駅��������é���I���u���딅�n�������,��������������ٖ��𘅽P   P   B���n������.���Π��S�������⚅���������М��\���&�����������1���������������P   P   &���p���������������՞��u���>���⚅�é����������������֔��Ȗ��ܘ��:�������e���P   P   ᙅ�͒��ԝ������a���𡅽[���u����������ߣ��b�������򑅽����E��������������$���P   P   И���������a���~�������𡅽՞��S�������"���-��������������虅�$���E���!���3���P   P   -�������7���K�����~���a�������Π��駅�e���E���$�������������/�������{���`���P   P   ����Л�����\���K���a�����������.���񜅽Y�������������y���Y�������ћ���������P   P   ]�������o������7�������ԝ���������񠅽���ԡ���������������������隅�o���ם��P   P   ȕ���������Л���������͒��p���n���ݜ��֠����������l�������%�������������������P   P   i����������̎�������������a���������������ܙ��.���7�������"�����Ì��=�������P   P   �������������������󗅽Ҋ������x���ҕ���������H��������������l�����������=���P   P   =���o���������������������ҍ��y�������E���֌��ˏ��j���n���*���������0�������P   P   Ì������ֈ��a�������튅�ߐ��W���1����������Ք��|���9�����������掅�.����������P   P   ��������������!��� ���������������I�������7�������j���x����������掅����l���P   P   "���u���z���ߍ��,���;�������%���>�������ѓ��3���ƍ��?���"�������������*������P   P   ���������������i���!���R��������������W�������쏅�|�������"���x�������n�������P   P   7���Ȟ������
������"�������ٛ��t������Փ��"���(�������|���?���j���9���j�������P   P   .���a�������ȏ��폅�����������������ޓ��ɒ�������(���쏅�ƍ������|���ˏ��H���P   P   ܙ��S���蘅�M�����������2����'������$��� �������"�������3���7���Ք��֌�����P   P   ����ᚅ�閅�w����@��������������E�������$���ɒ��֓��W���ѓ����������E�������P   P   ����斅�~���O���W���%���m���������������E������ޓ�������������I����������ҕ��P   P   ����m�����������"������ʧ��۞��Ý���������'�������t������>�������1���y���x���P   P   a�������q���{���5�������ܛ��$���۞���������������ٛ������%�������W���ҍ������P   P   ����H��������ƕ��񘅽Ψ��ܛ��ʧ��m�������2�����������R�����������ߐ�����Ҋ��P   P   ����ޕ��Q���`�����������񘅽�������%���@�����������"���!���;��� ���튅�����󗅽P   P   ������󔅽ɑ����������ƕ��5���"���W��������폅����i���,���!���������������P   P   ̎��׈��N������ɑ��`����{�������O���w���M���ȏ��
�������ߍ������a���������P   P   ��������ԍ��N���󔅽Q�������q�������~���閅�蘅������������z�������ֈ����������P   P   ����������׈�����ޕ��H�������m���斅�ᚅ�S���a���Ȟ������u�����������o�������P   P   @�����������φ��4���^���者�酅�}�������\��d����������������������
���`���.���P   P   .���情����ܑ���������[���҄������"���J����������T�����������ĉ��o�����������P   P   `�������ˉ��d����������c����������ߊ�������������􅅽w���؆������Q�����������P   P   
���猅�����\���Ƃ�����셅�w���������������؃��G�����������E���J���5���Q���o���P   P   ���-����������P����������􇅽t���h����������������������K���7���J�������ĉ��P   P   ������������5�������|�������w���@�������ˉ��内�J���p���@�������K���E���؆������P   P   �����������ڀ��N�������R�������������ڃ��h���=���]���7���@�����������w�������P   P   ��������G������6�������n���J������ˈ��\���$������L���]���p�����������􅅽T���P   P   ���������΍������@����������������������0����������=���J������G�����������P   P   d���C������������������܈������������������0���$���h���内�����؃���������P   P   \��������ʑ��ᑅ�ג��������������̂��s����������\���ڃ��ˉ�������������J���P   P   ��������L����������ډ���������݊��J���̂����������ˈ���������h�������ߊ��"���P   P   }����������Ќ��i������ˊ��t�������݊��������������������@���t��������������P   P   酅�j�������n���G���V���b���ń��t�����������������J�������w���􇅽w�������҄��P   P   者�F���Q���e�������	�������b���ˊ����������܈������n���R����������셅�c���[���P   P   ^���ف���������ጅ�f���	���V������ډ��ג�����@�����������|����������������P   P   4���y���싅� ���3���ጅ�����G���i������ᑅ���������6���N�������P���Ƃ����������P   P   φ������Ɉ����� ������e���n���Ќ������ʑ������΍�����ڀ��5������\���d���ܑ��P   P   ��������Ŏ��Ɉ��싅�����Q����������L�����������G�������������������ˉ�����P   P   ����q�����������y���ف��F���j��������������C������������������-���猅�����情�P   P   Dy���{��탅�ゅ�+}��ȃ��׉��M���҆������⋅�]���z���0���օ�����9��􇅽������P   P   ����w������	y�����p{��`���Y�������큅�u�������O���僅�]���D���C}��i~���x��n���P   P   ����s��C���%u��t~�������{���}��������W���	���o������׃��I}��H���~��������x��P   P   􇅽�~��
~��9���u|����������%|��5������΂��������.���р��?~���|������~���i~��P   P   9��6���Wr���|������'{��,{���������g}���~��-����~��-���T}��}��%����|��H���C}��P   P   ���X���E�������녅�ц��%����~���~��~���}��僅����~���섅��~��}��?~��I}��D���P   P   օ��M�������ņ��}�������4���'���聅�����~��̂�����􀅽G���섅�T}��р��׃��]���P   P   0��������~��o��������|��:�����������I���)���Ã���������􀅽~���-���.������僅�P   P   z���6���_���v������ۂ������T�������g����~��v���
��������������~�����o���O���P   P   ]���
���0���n����|��E|������r�������0������V���v���Ã��̂��僅�-������	�������P   P   ⋅������������E���U���t���恅�˃��������������~��)����~���}���~��΂��W���u���P   P   ����O�����������K���'�������㋅�����􌅽����0���g���I������~��g}��������큅�P   P   ҆��׃��-�������C���^�������B����������˃��������������聅��~������5����������P   P   M���󊅽����N���݌��<���T���Q���B���㋅�恅�r���T�������'����~�����%|���}��Y���P   P   ׉��򃅽~�������䃅�����ႅ�T�����������t�����������:���4���%���,{�������{��`���P   P   ȃ��B����y��}���
���X�������<���^���'���U���E|��ۂ���|������ц��'{����������p{��P   P   +}�����������������
���䃅�݌��C���K���E����|���������}���녅�����u|��t~�����P   P   ゅ�����}��M�������}�������N���������������n���v���o���ņ�������|��9���%u��	y��P   P   탅�&|���y���}�������y��~�������-�����������0���_����~������E���Wr��
~��C�������P   P   �{���u��&|���������B���򃅽󊅽׃��O������
���6�������M���X���6����~���s���w��P   P   �v���y��Sz��lw��~��Ys���r��\r���w��Bx��bu���z���v��Ou��dw���s���y��&y��v��_|��P   P   _|��8����{��v������z��Mr��Sv��ty���{���u���q��A}���v��Gu���r��K{���z���{��S}��P   P   v��	z��Pv���w���y��"o��m}��&}��rx��Dr���w��{t���t��Nv��v���|��W|��Hu���u���{��P   P   &y���|��|��x��s����l���t���}��x���y��v��3~��"{��Zz��xv���y���z���r��Hu���z��P   P   �y��w�������x��}w��P}��m{��I���r��|��w{���w���u��Ey���|��Jz��oz���z��W|��K{��P   P   �s��`r��[u���{���n���t���u���|��Gx���z��{���s��yu��Bv���r���z��Jz���y���|���r��P   P   dw��}���|���{���x��}��ct���s���v���w��G|��,t���s��|���q���r���|��xv��v��Gu��P   P   Ou��Xu���t���w���r��#y���v��{t��y���t��Oz��Wy��u��lz��|��Bv��Ey��Zz��Nv���v��P   P   �v���r���v���x��8|��\{��bv��<q���x��x��;y��Cy���t��u���s��yu���u��"{���t��A}��P   P   �z���q��[|��Y{�����e���f~���x���v���v���s���v��Cy��Wy��,t���s���w��3~��{t���q��P   P   bu���q��z���x��y��@|��u���x���v���s��st���s��;y��Oz��G|��{��w{��v���w���u��P   P   Bx��"o���w�����Nx���}��~���x��W����v���s���v��x���t���w���z��|���y��Dr���{��P   P   �w��Av��z��@}���{��mv��]|���w���|��W����v���v���x��y���v��Gx���r��x��rx��ty��P   P   \r���n���{���z���v���x���p���p���w���x���x���x��<q��{t���s���|��I���}��&}��Sv��P   P   �r��y��7t��Q}���w�� ~��|���p��]|��~��u��f~��bv���v��ct���u��m{���t��m}��Mr��P   P   Ys��e~��z|��5y������}�� ~���x��mv���}��@|��e���\{��#y��}���t��P}���l��"o���z��P   P   ~�� q��Qs��x��{w������w���v���{��Nx��y�����8|���r���x���n��}w��s����y�����P   P   lw��{x���y���}��x��5y��Q}���z��@}������x��Y{���x���w���{���{���x��x���w��v��P   P   Sz���z��J����y��Qs��z|��7t���{��z���w��z��[|���v���t���|��[u������|��Pv���{��P   P   �y���~���z��{x�� q��e~��y���n��Av��"o���q���q���r��Xu��}��`r��w���|��	z��8���P   P   �l��gk���k���i���p���t���p��by��	q��uv��zu��9u���v��u���t���q���u��g���n���h��P   P   �h��Np���g��eu��jj���q���s���u��[q��p���w���q���r���p��it���p���r��l���s��Fj��P   P   �n���u���h���w��Qv��on��Ss��l���q��"s��_p��?x���u���q���s���p���o��	r���r���s��P   P   g��6k��kk���g���j���n���v���l���o��t��o��o���o���j�� r��Ko��Xo��bq��	r��l��P   P   �u��Pq��Aq��.t���o��!r���t��Bi���p���o���l���n���n���l���n��4o���m��Xo���o���r��P   P   �q��Ts���n���l���u��ws���r��Xl��wq��r��Hl��	u���t���x���s���n��4o��Ko���p���p��P   P   �t��On��ws���m��	q���s��p��hu��kt���r��fk���s���s���j��Jr���s���n�� r���s��it��P   P   u���w��?x���v��Fu���y���t���x��p���o���m��zm���u���m���j���x���l���j���q���p��P   P   �v��s��gt���p���m��#r���n���t��Cu���q���v���o�� r���u���s���t���n���o���u���r��P   P   9u��ez��0s���r��Vq���p���r��Nv��9y��5x���s���q���o��zm���s��	u���n��o��?x���q��P   P   zu���x���w��!t���r���q��Hp���w���v��Fv���w���s���v���m��fk��Hl���l��o��_p���w��P   P   uv��w���p��p��r��p��kt���p���q���n��Fv��5x���q���o���r��r���o��t��"s��p��P   P   	q��,{���w��#p���t��x��y���x��p���q���v��9y��Cu��p��kt��wq���p���o���q��[q��P   P   by���y��~s���u���q���v���y���v���x���p���w��Nv���t���x��hu��Xl��Bi���l��l���u��P   P   �p��Ft��Pn���n��Et���q���x���y��y��kt��Hp���r���n���t��p���r���t���v��Ss���s��P   P   �t���p��Gy��<w��o���q���q���v��x��p���q���p��#r���y���s��ws��!r���n��on���q��P   P   �p��Jt���o��s��Kp��o��Et���q���t��r���r��Vq���m��Fu��	q���u���o���j��Qv��jj��P   P   �i���o���s���l��s��<w���n���u��#p��p��!t���r���p���v���m���l��.t���g���w��eu��P   P   �k���l��n���s���o��Gy��Pn��~s���w���p���w��0s��gt��?x��ws���n��Aq��kk���h���g��P   P   gk��Ns���l���o��Jt���p��Ft���y��,{��w���x��ez��s���w��On��Ts��Pq��6k���u��Np��P   P   mq��^m���n��Ts���d���h��g���e��a���a��Ze��A_���f��7d���g��i��ff��^p��r���j��P   P   �j���e��Di���e��Ke��ne��j��&h��e��i���d���f���b���e��g���j���c��af��f��i��P   P   r��*g���p���h���a���p��`���f��'d��1n���c��rb��Gi�� i���h���d��e���j���f��f��P   P   ^p��rh��bj���t��'`���o���i���g��/l���d��n��g��i���j���j��ve���i��?k���j��af��P   P   ff���k��!`��uh�� j���d��Id��3f���q���d��Ih���k���h��"j���j���h���l���i��e���c��P   P   i��rj���n���h��2l���h��dg���e��(i���d��6j��'h���a���d���f��5e���h��ve���d���j��P   P   �g���a��Ed���j���f��}^���g���i���h��Qf��l��<h��|d���h���e���f���j���j���h��g��P   P   7d��.e��+d��qf��wj��Bb���f���e���c���j��>j��Zj��na��l���h���d��"j���j�� i���e��P   P   �f���g���i��^i��xj���g���j���j��a�� h��Gf��=h��hj��na��|d���a���h��i��Gi���b��P   P   A_���b��Gb���h���g��wi���f��Cd��1_���`��f���c��=h��Zj��<h��'h���k��g��rb���f��P   P   Ze��f��Oc��Wi���m��Dl��7p��if��Rc��Cg��hc��f��Gf��>j��l��6j��Ih��n���c���d��P   P   �a��Yh���k���g��7n��gf��h��]l���h��Fo��Cg���`�� h���j��Qf���d���d���d��1n��i��P   P   a��S^���a���j���j���g��a��^g��k���h��Rc��1_��a���c���h��(i���q��/l��'d��e��P   P   �e���l���b��h���m��Vd��Vh���e��^g��]l��if��Cd���j���e���i���e��3f���g���f��&h��P   P   g��Jb��j���j��gn���g��c��Vh��a��h��7p���f���j���f���g��dg��Id���i��`��j��P   P   �h���c��`���i���h��2j���g��Vd���g��gf��Dl��wi���g��Bb��}^���h���d���o���p��ne��P   P   �d��_j���k��jg���h���h��gn���m���j��7n���m���g��xj��wj���f��2l�� j��'`���a��Ke��P   P   Ts��Bk���f���k��jg���i���j��h���j���g��Wi���h��^i��qf���j���h��uh���t���h���e��P   P   �n���k���a���f���k��`��j���b���a���k��Oc��Gb���i��+d��Ed���n��!`��bj���p��Di��P   P   ^m��_c���k��Bk��_j���c��Jb���l��S^��Yh��f���b���g��.e���a��rj���k��rh��*g���e��P   P   Z���^��[���Z��.^��z^��<b��C^��*j��h��tc���i���f��|a��1`���a��.Z���^��=X��Za��P   P   Za��{[��Ic��m[��qh��Je���^��;_��d���g���b��#j��
f���e��u^��a���b���g���[��6^��P   P   =X��^W��[��![���_���\���`��_j���`���[��z`���a���\��^��1a���e��~c���]���a���[��P   P   �^��Ja���b��Z��qi��^���W��c���^��M^���[��d���`��^^��][��	`���`���Y���]���g��P   P   .Z��Z��Bh���W���\��-e��W_��ug��*W���b��b���\��'b���_�� `��`��`���`��~c���b��P   P   �a���[��2_���b���\��)_��8`���h��*`��,]���d��Z\��b���]��`��Nb��`��	`���e��a��P   P   1`���l���c��"_���e��!h���e���]���\�� ^���b���[��c���d��Oa��`�� `��][��1a��u^��P   P   |a��Zb���d��E^���]��c��5d��!\���d���a��E_���^��w`���d���d���]���_��^^��^���e��P   P   �f��c���`��ac���e��ub���d���_���k��}f��cZ��`���a��w`��c��b��'b���`���\��
f��P   P   �i��f���h���a���`���`��b���f��j���g��e���h��`���^���[��Z\���\��d���a��#j��P   P   tc��`���f���b��!\��_��e]���a��0e���b���c��e��cZ��E_���b���d��b���[��z`���b��P   P   h��Ec��c���a��>]��3g��lb��u^���a���`���b���g��}f���a�� ^��,]���b��M^���[���g��P   P   *j��jh���f��Kc���^���c��i���b���b���a��0e��j���k���d���\��*`��*W���^���`��d��P   P   C^���^���g���`��o^��5c���c���e���b��u^���a���f���_��!\���]���h��ug��c��_j��;_��P   P   <b��:f���d���b���Y���f���h���c��i��lb��e]��b���d��5d���e��8`��W_���W���`���^��P   P   z^��-j���c��x_��^b��Ba���f��5c���c��3g��_���`��ub��c��!h��)_��-e��^���\��Je��P   P   .^��S[���b���`���d��^b���Y��o^���^��>]��!\���`���e���]���e���\���\��qi���_��qh��P   P   �Z��^���^��=`���`��x_���b���`��Kc���a���b���a��ac��E^��"_���b���W��Z��![��m[��P   P   [��^���h���^���b���c���d���g���f��c���f���h���`���d���c��2_��Bh���b��[��Ic��P   P   �^���W��^��^��S[��-j��:f���^��jh��Ec��`��f��c��Zb���l���[��Z��Ja��^W��{[��P   P   wP���X���Y��S���[���X��KX���[���R��{P��S��|S��5L���\���U��W��h_���V���W��F[��P   P   F[���_���Z���]��,V��&V���R���V��)W���K���R���P���O��TU���W���R��cV���T���]���\��P   P   �W���a��`X��EZ���[���Q��9]��NP���Z���V���]��SY��;W���[��mV��jU���X��?V��1U���]��P   P   �V���V���Y��uS���X��T���`��AV���Q���_��|X���V��U���]��)Z��QZ��NT���]��?V���T��P   P   h_���[��UX��O^��!]���U��=W���T��T���\��&V���U��nU��mV��V��hX���S��NT���X��cV��P   P   W��S[���R���T���[��T���T���R��)Y���^��dP��:Z���]��Y��JY���V��hX��QZ��jU���R��P   P   �U��_P��xX���W���U���S���W���X��-U���[���R���Y��'Z���M���[��JY��V��)Z��mV���W��P   P   �\���U���T���Z��eX��~U��=V��rY��Y��LZ���Z��bW���]���G���M��Y��mV���]���[��TU��P   P   5L��JT���T���T���T��uV���S���P��S���L��3W��jV��U���]��'Z���]��nU��U��;W���O��P   P   |S��5S���S��RX���Y��gW���W��xS���R���N���Q���\��jV��bW���Y��:Z���U���V��SY���P��P   P   S��gX��U���V���Z��;Z��YZ���Z���V���T��Y���Q��3W���Z���R��dP��&V��|X���]���R��P   P   {P��DU��;R���Y���X��kW���V���Y���W��RR���T���N���L��LZ���[���^���\���_���V���K��P   P   �R��PU���S���U��C\��W��U��mW���X���W���V���R��S��Y��-U��)Y��T���Q���Z��)W��P   P   �[��vN���T��sZ��[��MZ���S���U��mW���Y���Z��xS���P��rY���X���R���T��AV��NP���V��P   P   KX��W��T���W��IZ��AT��0S���S��U���V��YZ���W���S��=V���W���T��=W���`��9]���R��P   P   �X��vP���V��cT��vY��Z��AT��MZ��W��kW��;Z��gW��uV��~U���S��T���U��T���Q��&V��P   P   �[���[��S���Y��W��vY��IZ��[��C\���X���Z���Y���T��eX���U���[��!]���X���[��,V��P   P   S���Z���Y��TV���Y��cT���W��sZ���U���Y���V��RX���T���Z���W���T��O^��uS��EZ���]��P   P   �Y��MY��UT���Y��S���V��T���T���S��;R��U���S���T���T��xX���R��UX���Y��`X���Z��P   P   �X���f��MY���Z���[��vP��W��vN��PU��DU��gX��5S��JT���U��_P��S[���[���V���a���_��P   P   �V��yL���K��)V��jK��S��$Q��$P���T��X��U��XV��oV��!O���S��QQ��_L���O���Q���G��P   P   �G���M���D��<N���K���M��V��NP���O���U��OX���Q��	Y���P��7R���U���N���I���N���F��P   P   �Q���J��N��1P��bN��R���M���O��VQ��_P��Q��uM���R��O���K��UO���L���S���P���N��P   P   �O��L��'J��VV��*F��	S��iQ���P���T���H��O��+K��|P��AL���K��IT���P���Q���S���I��P   P   _L��vQ��I��	P���L��)O���R��~H��yZ��{I���N��PT��R���R���N���O��Q���P���L���N��P   P   QQ��-O��FT��O���O���R��V���P��FQ��O��O��tP���G���L���K���Q���O��IT��UO���U��P   P   �S��NL���O���S��qO���M��}M��cR���Q���G��P���R���J���Z��nO���K���N���K���K��7R��P   P   !O���R���S��P��S���Q��S��QP��7M���N���N��pQ���J��\���Z���L���R��AL��O���P��P   P   oV���U���V��+Q���N���S��"V���Z���S���X��QU��P���L���J���J���G��R��|P���R��	Y��P   P   XV���V���P���Q���P��OQ��uP���Q�� T��pW��}T���G��P��pQ���R��tP��PT��+K��uM���Q��P   P   U���S��
O���O���Q���N���Q��RL��R��ES��%V��}T��QU���N��P��O���N��O��Q��OX��P   P   X��nT���V���S���R��XN���P��/Q��]P���X��ES��pW���X���N���G��O��{I���H��_P���U��P   P   �T���S��HQ���O��L���O��]P��`Q��O��]P��R�� T���S��7M���Q��FQ��yZ���T��VQ���O��P   P   $P���X��R��wP��O���P���V���T��`Q��/Q��RL���Q���Z��QP��cR���P��~H���P���O��NP��P   P   $Q��'P��
W���O���S���O�� S���V��]P���P���Q��uP��"V��S��}M��V���R��iQ���M��V��P   P   S��	K��NU��yR���N���P���O���P���O��XN���N��OQ���S���Q���M���R��)O��	S��R���M��P   P   jK��{P��DS���Q��dN���N���S��O��L���R���Q���P���N��S��qO���O���L��*F��bN���K��P   P   )V��<P���P���O���Q��yR���O��wP���O���S���O���Q��+Q��P���S��O��	P��VV��1P��<N��P   P   �K���N���D���P��DS��NU��
W��R��HQ���V��
O���P���V���S���O��FT��I��'J��N���D��P   P   yL���G���N��<P��{P��	K��'P���X���S��nT���S���V���U���R��NL��-O��vQ��L���J���M��P   P   TJ��'M���L��;G���C��F��KF���A���B���?��	B��?���D��??��C���E���D���G��]L��GL��P   P   GL��AF��P��#D��L���K���E���D��LF��eE��eA���C��fB��ZH���E��/E���K��:O��eD��L��P   P   ]L��nF���H��J��)G���J��ZA���I��PF��4H��1A��VH���E��E��uJ��G��D���D��'I��eD��P   P   �G��fM���J���I��1K���G���>��4F��5G���F���H���G���I��'B���K���E��sI��>?���D��:O��P   P   �D���C��nN���B��,C���I��'E��I���C���D��IM��)G��cJ��5G��7K���C��2A��sI��D���K��P   P   �E��qD��	H��oJ��
D���J���?���H���E���@���M��?F���E���G���J��J���C���E��G��/E��P   P   C���P���D���A��9H���N���E��9D��!M��BJ��NN��E��>D�� C���?���J��7K���K��uJ���E��P   P   ??��DD���H���B���C���E���C��;E���C��LD�� D��4D��qE���J�� C���G��5G��'B��E��ZH��P   P   �D��UA���>���F��bJ���C���>��3@��[B���E�� D��RJ��_P��qE��>D���E��cJ���I���E��fB��P   P   ?��D���H���D��}G��G��)G���G���B���B��^C��fD��RJ��4D��E��?F��)G���G��VH���C��P   P   	B��
>��/F��&H��ZC���D��yE��}H���F��w@���<��^C�� D�� D��NN���M��IM���H��1A��eA��P   P   �?���@���F���D���F���K��vI��nG��1F��ND��w@���B���E��LD��BJ���@���D���F��4H��eE��P   P   �B��u@���H���H���F��?J��AI��_F��nH��1F���F���B��[B���C��!M���E���C��5G��PF��LF��P   P   �A��E���E��0F���G���G��B��HC��_F��nG��}H���G��3@��;E��9D���H��I��4F���I���D��P   P   KF���D���?���D��D��
K���E��B��AI��vI��yE��)G���>���C���E���?��'E���>��ZA���E��P   P   F��GN��4C���E���H��.D��
K���G��?J���K���D��G���C���E���N���J���I���G���J���K��P   P   �C��]C��I��WB���K���H��D���G���F���F��ZC��}G��bJ���C��9H��
D��,C��1K��)G��L��P   P   ;G���E���G��	B��WB���E���D��0F���H���D��&H���D���F���B���A��oJ���B���I��J��#D��P   P   �L���J��*R���G��I��4C���?���E���H���F��/F���H���>���H���D��	H��nN���J���H��P��P   P   'M���A���J���E��]C��GN���D��E��u@���@��
>��D��UA��DD���P��qD���C��fM��nF��AF��P   P   2��v9��8?��Q9��4H���;���?���E���B���D���J���F���A�� J���>���;���C��i<��r5���>��P   P   �>��(<���?���:���=��{<��|:���B��B���@���?���C��7=��	@���B��>��<��e=���>��B@��P   P   r5��A���;���9���=���;���E���@��<��+@���B��C���A��>A��D<��>��VE���<���:���>��P   P   i<��P:��>���7���A���9���E��c@���9���B��)?���A���<���C���A���9���@���F���<��e=��P   P   �C��1?���9��,B��D���>��NA��iH��>��I���8��7���7���7���;��eC��xE���@��VE��<��P   P   �;���D���;���?��W?��=��>���<��8;��l@���6��z<��"J��D���>���4��eC���9��>��>��P   P   �>���;��`?��7C���<��9���A��B���9���D��K=���=���I���9���E���>���;���A��D<���B��P   P    J��'D��;��G��_C���B���@��^I���B���@���@���8���C���3���9��D���7���C��>A��	@��P   P   �A���E��XA���A���=��/A��}E��_A��lC��4=��B���:���=���C���I��"J���7���<���A��7=��P   P   �F��@���@��fC��j@��E?���B���A���B��~C��TC���G���:���8���=��z<��7���A��C���C��P   P   �J���H���B��eA��@A��D��I?��E@��F?��J��fH��TC��B���@��K=���6���8��)?���B���?��P   P   �D���F��7>��$>���>��=���<���?��?@��=>��J��~C��4=���@���D��l@��I���B��+@���@��P   P   �B���D��^?���>��E���<��$<���>��B��?@��F?���B��lC���B���9��8;��>���9��<��B��P   P   �E��B��YB���?��e@��p>���A���E���>���?��E@���A��_A��^I��B���<��iH��c@���@���B��P   P   �?���C��B��IF��d@���=��$>���A��$<���<��I?���B��}E���@���A��>��NA���E���E��|:��P   P   �;��I>���=���B��?��pA���=��p>���<��=��D��E?��/A���B��9��=���>���9���;��{<��P   P   4H��A���=��E���;��?��d@��e@��E���>��@A��j@���=��_C���<��W?��D���A���=���=��P   P   Q9���=��<���E��E���B��IF���?���>��$>��eA��fC���A��G��7C���?��,B���7���9���:��P   P   8?��?:��>=��<���=���=��B��YB��^?��7>���B���@��XA��;��`?���;���9��>���;���?��P   P   v9��KA��?:���=��A��I>���C��B���D���F���H��@���E��'D���;���D��1?��P:��A��(<��P   P   E��9���5��1:���5���9���6���/���1��&3���'��3���3���,���7��;���1��o<��t5��f6��P   P   f6��<���1��]>���4���1��4:��V4��2���6��>5���2��f:���1���2���:���4���2��t=��x6��P   P   t5��a9���:���:��w>���5���8��&7��F9���2���4���.��r2��|5��9���9���2��:;��X9��t=��P   P   o<���;���7���7���5��_7��03���-���6��
3��S5��h9��7���7���-���8�� .���1��:;���2��P   P   �1��":��h3���9��K4��3���4���-���7���6��68��@��b9��H?��8��%7��[8�� .���2���4��P   P   ;��%6��(7���6���8���5���?���6��:��(7���7��n9��@-��0��36���;��%7���8���9���:��P   P   �7���3��H6���5��C5��/8��I5���4���5���0���5���:��R0��D;���6��36��8���-��9���2��P   P   �,���4��5��U5��L1���7��*3���)��U4��z5��P7���>���2��x9��D;��0��H?���7��|5���1��P   P   �3���1��:��5��E0��4��v5��b5���3��h7��Q5��S7���5���2��R0��@-��b9��7��r2��f:��P   P   3���1��6/��A4��2���8���0��2���3��2���0���/��S7���>���:��n9��@��h9���.���2��P   P   �'��/��7���3��65��6��5��S4��t4���-���-���0��Q5��P7���5���7��68��S5���4��>5��P   P   &3���-��6��O7���7���7���8��8��|8��V5���-��2��h7��z5���0��(7���6��
3���2���6��P   P   �1��w5���5���6��r5���6���7���7���0��|8��t4���3���3��U4���5��:���7���6��F9��2��P   P   �/��1���1���5���4���4��9���5���7��8��S4��2��b5���)���4���6���-���-��&7��V4��P   P   �6���4��.6��S0��=6��6��N<��9���7���8��5���0��v5��*3��I5���?���4��03���8��4:��P   P   �9��^3��b8���5��"4���:��6���4���6���7��6���8��4���7��/8���5��3��_7���5���1��P   P   �5���6��q4���3��a0��"4��=6���4��r5���7��65��2��E0��L1��C5���8��K4���5��v>���4��P   P   1:��>7���7���5���3���5��S0���5���6��O7���3��A4��5��U5���5���6���9���7���:��]>��P   P   �5��X9���7���7��q4��b8��.6���1���5��6��7��6/��:��5��H6��(7��h3���7���:���1��P   P   9��h;��X9��>7���6��^3���4��1��w5���-��/���1���1���4���3��%6��":���;��a9��<��P   P   &)��^,��,���.���(��F0��+0��A5���2��91���6���.���3��3��X0��_/���+��U+���0���*��P   P   �*�� '��.��'+��6-���2��=-��e*��c3���-�� 7��%5��p-��3��'-���(��n4��x1��&��1��P   P   �0��<(���.��*��8$��j1���+��?*���2���2���.��)4���0��A0��3��-��A+���.��v'��&��P   P   U+��(.��Q)���0���+���2���1���5���4��f.��C-���'��.-���*���0��I3��(8���0���.��x1��P   P   �+��&*���0��>+��I.��`0��I/���0��:1���#��//���,���0��L-���-���(��](��(8��A+��n4��P   P   _/���)��Y2��v.���*��Q,���)��c+��83���+���2��/���+���.���+���3���(��I3��-���(��P   P   X0���2���/���+���0��4���/��[-���5���-��g-��d+���(��x2��D)���+���-���0��3��'-��P   P   3��h.���1��3.��%2���+���1���3��U3��.��C,��r,��-���8��x2���.��L-���*��A0��3��P   P   �3��Z2���-��/��K7��#1���*���5���/���/���.��|0���+��-���(���+���0��.-���0��p-��P   P   �.���6��D3��a1��+2��>5���1���2��u0���3���5���/��|0��r,��d+��/���,���'��)4��%5��P   P   �6���4��%1��#1���0��L*���-��23���2��\3���7���5���.��C,��g-���2��//��C-���.�� 7��P   P   91���6��51���,���.���.��i-��*0��W-��(3��\3���3���/��.���-���+���#��f.���2���-��P   P   �2���0���0��/.���,��L1��|/���0��+��W-���2��u0���/��U3���5��83��:1���4���2��c3��P   P   A5��#4���2��j3���1��h/��(��~%���0��*0��23���2���5���3��[-��c+���0���5��?*��e*��P   P   +0��V.��0���.���/��.���-��(��|/��i-���-���1���*���1���/���)��I/���1���+��=-��P   P   F0��/��c/���/��P3���)��.��h/��L1���.��L*��>5��#1���+��4��Q,��`0���2��j1���2��P   P   �(��,��=4��.-��,;��P3���/���1���,���.���0��+2��K7��%2���0���*��I.���+��8$��6-��P   P   �.��Q+��0���*��.-���/���.��j3��/.���,��#1��a1��/��3.���+��v.��>+���0��*��'+��P   P   ,���,���.��0��=4��c/��0���2���0��51��%1��D3���-���1���/��Y2���0��Q)���.��.��P   P   ^,���)���,��Q+��,��/��V.��#4���0���6���4���6��Z2��h.���2���)��&*��(.��<(�� '��P   P   +%���)��D'��~&���)���!���$���#��
$��N!���$���"�����A(���#��� ��-��Y$��f'��#+��P   P   #+��=)��-��M'��	*��='��m'���(���"��� ��������G ��V#���*���(��0#��*���(��T'��P   P   f'��:,��'��s'���(���$���!��'������"��o'��a%��B'���#�����"��S)������-���(��P   P   Y$���$���&���$��2)��e"��� ���&��8"���'��+��D'���'���'��4,��H ��*#��%�����*��P   P   -��o&���'���'��(+��'&���&���&��i���*���%��G��Y%��5���$��7,���"��*#��S)��0#��P   P   � ���)��(%��m%���$��]'��o&���&����G*��7&���#���1��$-���(��d!��7,��H ���"���(��P   P   �#��-#���$���#���&��� ���$���%�����1)���&���$��{-������)���(���$��4,�����*��P   P   A(���"��:&���#��)��	#���!��u(��)"���#���)��D#���,��������$-��5���'���#��V#��P   P   ���F"���"��2#��C���!���(��� �� ��� ��T&���$��*&���,��{-���1��Y%���'��B'��G ��P   P   �"��  ��_$���#��O"������&���!��� ���#�����9$���$��D#���$���#��G��D'��a%�����P   P   �$��E �����1$���%���*���%��8!��2 ��/$�������T&���)���&��7&���%��+��o'�����P   P   N!���#��[!��C*���"���#���$��%��W$��!��/$���#��� ���#��1)��G*���*���'���"��� ��P   P   
$��u��A��%��B(��r$���&���$��u,��W$��2 ��� �� ��)"�������i��8"������"��P   P   �#��� ���$��u ��A#��_&��H.��.0���$��%��8!���!��� ��u(���%���&���&���&��'���(��P   P   �$���"���&��w'�� &���'��P%��H.���&���$���%���&���(���!���$��o&���&��� ���!��m'��P   P   �!���#���#���������$���'��_&��r$���#���*������!��	#��� ��]'��'&��e"���$��='��P   P   �)�� '���'��0&��� ����� &��A#��B(���"���%��O"��C��)���&���$��(+��2)���(��	*��P   P   ~&���*���"��2%��0&�����w'��u ��%��C*��1$���#��3#���#���#��m%���'���$��s'��M'��P   P   D'��G&��'$���"���'���#���&���$��A��[!�����_$���"��:&���$��(%���'���&��'��-��P   P   �)��4)��G&���*�� '���#���"��� ��u���#��E ��  ��F"���"��-#���)��o&���$��:,��=)��P   P   !��J��R����������S��0���"��$��?���'�����?��,�������l�������P   P   ���������P���������� ��� ��g(���$���"���(��b"������ ����������i��P   P   ��D��������"������!��q"���"����������������(#���"��K!��m!��L ����P   P   l��������~��������������v��������� ��o�����<��#��������m!�����P   P   ���A�����4�����$��0�� ��r��i"�����j!����V"��������%�����K!�����P   P   ����x�����d��m ��p��y$��� ����U����������5��������#���"��� ��P   P   ,��������f ��y���!�����;��� ��j��T��b������"����5����<��(#�����P   P   ?���"����~�����# ��$��P��~!��Z ��\��!���������"�����V"��������b"��P   P   ���� ��d!��
$��$��� ���#�����"���#��������������������o������(��P   P   �'��}#���!��A��#��� ���������%��f%���#��c����!��b����j!��� ������"��P   P   ?�����$��i��E��t!���!�����&��	 ��!���#�����\��T��U�����������$��P   P   $��>��p#��s����� ��L������!�����	 ��f%���#��Z ��j����i"��������g(��P   P   �"���$���'��� ��D��/�����������!��&���%��"��~!��� ��� ��r��v���"��� ��P   P   0��'���������������������������������P��;��y$�� �����q"��� ��P   P   S���#�����E�����T��A��������L���!������#��$�����p��0������!����P   P   ���!������!��<#��d!��T�����/�� ��t!��� ��� ��# ���!��m ��$�����������P   P   ���������\ ��!��<#�������D�����E��#��$�����y��d���������"����P   P   ���>�����!��\ ���!��E������ ��s��i��A��
$��~��f �����4��~�����P��P   P   R�����n�����������������'��p#��$���!��d!�������x�������������P   P   J��������>������!���#��'���$��>�����}#��� ���"�������A�����D�����P   P   z�������&��������h�����,��3��O��5	�����o����������~��������P   P   ������)��/��h��%�����A��]���
�����G���
��������d�������������P   P   ������F��������B�����:�������������[�������e������������P   P   ~��l����#��'�����C�������������)��K��z�����������d�������P   P   �����N������������J��,��!�����,����I��������������������P   P   ��������������������y��x�������������f�����7��������e��d��P   P   �����������������i���������������������������������������P   P   o��������������J��a�������i��y��������������f��I��z�������P   P   ���B�������a��'��.����������������@������������K��[���
��P   P   5	��D�������T����������� ��~�����z��������������,��)����G��P   P   O��������x��q��p	������������e��������y������������������P   P   3��������
��?��1�����:����?����~�����i�������!���������
��P   P   ,��Z��������L����� ������������� �����������x��,��������]��P   P   ��������������������S�����:���������������y��J�����:��A��P   P   h��l��������`��
�������� ����������.��a��i������C��������P   P   ���������%��������
��������1��p	�����'��J�������������B��%��P   P   ������@��P�������`�����L��?��q��T��a��������������'�����h��P   P   &����������P��%������������
��x������������������#�����/��P   P   �����������@���������������������������������N����F��)��P   P   �����������������l����Z��������D��B��������������l��������P   P    ��8����������������1��-��B��������h�����������d�������d	��P   P   d	���	��V���
������	��������������<��]�����/
��E������
�����	�����P   P   ������	���
����<��:�������;�����%�����������^�����������	��P   P   �����������=������
�������V����'��:��>�����Z	��1��w
�������P   P   d�����D����������������%����x
�����5��#����|�����1������
��P   P   ��������?
�������������������������v�����V	�����|��Z	��^�����P   P   ���B��v��@��������\�����!��x��P�����w
��/ ����V	����������E��P   P   ���J����/��1��}��_	���
��J��������������	��/ �����#��>�����/
��P   P   h��]��%������	��I����������������:��������w
��v��5��:��������P   P   ���������������^�����������������:��������������'��%��]��P   P   ���7��c�������������F������������������P����x
�������<��P   P   B��)��������
��*��]���������������������x�������V��;�����P   P   -���������������������&������������J��!�����%�����������P   P   1������������
�����
����������F���������
������������������P   P   ��������W������������
�����]���������_	��\���������
��:�����P   P   ������]��������V����������*�����^��I��}�������������<���	��P   P   ��������������������
�����
���������	��1�����������=�������P   P   ���u�����;�������W��������������������/��@��?
���������
���
��P   P   ��������������]�������������c�����%����v����D������	��V��P   P   8�������u����������������)��7�����]��J��B��������������	��P   P   ������	��N������w��J���������������������@ ��"�������� ��2��l	��P   P   l	��p��!��5��r������ ��� ��������� ��&��#��K��W�����U��a��W��g��P   P   2��<�����������a��S�������e���*�������Y�������U��� �����2��	��W��P   P    ��������s��!�����F��=��g��(��v��4
�����^��c�����^������2��a��P   P   ������t�����O��|��������r���"��*�����D�����<��������^������U��P   P   ���������:�����o��7��� ��������������������
������������� �����P   P   "������������ ��������� �������/��L������������
��<��c��U��W��P   P   @ �����^ ��Q��������������I������G�����, ��o����������^������K��P   P   ����(�����k���S��V���#��(���R��� �����������, ��������D�����Y���#��P   P   ���� ��*���������z���9 ����n�����r�����������L��������4
������&��P   P   ��������8������� ��	��0���M �����m�������r������G��/�����*��v��*���� ��P   P   �������@���t���u��N��y���������V ��m������� ������������"��(��e������P   P   ��������������������:���	��{���������n��R��I�������r���g��������P   P   J����������L ��^���	���
��
���	�����M ����(������ �� �����=����� ��P   P   w���
��`����������l��^���
��:��y��0���9 ��#��������7������F��S��� ��P   P   ��T��)��������������l���	�����N��	��z���V����������o��|�����a�����P   P   ��*���������R����������^����u��� �����S������ �����O��!�����r��P   P   N�����V��A�������������L ������t�����������k���Q�����:�����s�����5��P   P   �	��E��[���V������)���`��������@���8��*�����^ ���������t��������!��P   P   ����E�����*��T���
������������������� ��(����������������<��p��P   P   ;���q􄽄���<���������������������������������������g�������J�������X�������P   P   ��������(����������������������g��u������o��
������'�������Z������#������P   P   X�����`���j���������������������� ��s���� ������>��<��4�������������#���P   P   �������X���(���b������������������G�����������+�������������J��������������P   P   J������������������������������ ��N���������<������P����������J�������Z���P   P   ����>������������������3�������m���]�������7���������s�������������4�������P   P   g���������h������S���#������B������A���	�����4�������s���P�������<��'���P   P   ������+�������b�������V �� ����������������������4������������>�����P   P   �����������v���m��S �������������@���i���Y��� �������������<���+�������
���P   P   ���
 ���������%������c������ ��S����������Y�����	���7���������� ��o��P   P   ������7�������������]��j������ ��������i�������A���������������s������P   P   ���������n������1������������������ ��S���@����������]���N���G���� ��u���P   P   ����^��������o���L���H������������������� ��������B��m���� ��������g��P   P   �����������������������󄽚�������j��������� �������������������������P   P   �����������������5���K�����H������]��c������V ��#���3������������������P   P   ������������ ��*������5�������L���1�����������S ������S����������������������P   P   ��������������n���*�������o���������%��m��b���������������b�����������P   P   <������������������ �����������n���������v�������h���������(���j������P   P   ��������{���������������������������7����������+��������������X���`���(���P   P   q�������������������������^��������
 ������������>����������󄽤���P   P   ������������s� �-���{򄽫�����턽�����3y�$���2�y�������P   P   �������O����H���-������鄽���h턽�鄽�s섽_�����G�������:�������P   P   �������X�����Y���J�C�n�tꄽ�󄽩���b����������넽9����u􄽎���:���P   P   y�_�������j���������
����Q�
󄽽넽g����/�	�������u􄽆���P   P   2�������������l��턽 �����)�d񄽎��������鄽�����G���P   P   $����􄽢�B턽Z���p����������������]������i���d�������������	�9�������P   P   y�.����� ꄽ���������񄽽􄽸넽���������!������������/󄽊넽_�P   P   3W턽m���^5�I����섽H�n鄽q��� 넽���L�����d������������s섽P   P   ��������󄽿섽������􄽛�^����u����!�i�������g�����P   P   ������򄽘ꄽ�턽�섽V����N넽� 넽�������d񄽽넽b񄽭鄽P   P   �턽����鄽>턽�鄽Q����񄽾ꄽ�턽�넽��N넽^������]���)�
󄽩���h턽P   P   ���턽�ꄽ���D���������섽���넽󄽛�q��������Q������P   P   �􄽇��鄽����������������6� ������턽����n鄽�넽�������tꄽ�鄽P   P   {�H򄽇����섽~턽���X �����6��섽�ꄽV񄽊�H񄽽������
���n򄽥�P   P   -���脽����"������q���X �������������섽��섽����� ���C����P   P    ������� �V턽�����������������Q����턽��I�������p����턽����J�-P   P   s������������焽V턽�~턽����D�鄽�ꄽ�섽5񄽶���Z���l�j���Y���H���P   P   ��@�������]儽�� �"����섽�������>턽���^ ꄽB턽�������������P   P   ����v���������������������������鄽�ꄽ鄽��m���������������X�O�P   P   ��������v���@���������脽H򄽇�턽����������W턽.�������_�����������P   P   �����鄽}脽�섽�ꄽ�섽x)ꄽ��U􄽉(넽X����섽�ꄽ�턽�焽�섽鄽P   P   鄽焽ꄽ�ꄽ�鄽\턽}脽N턽8�O~ꄽ������"鄽�넽
턽�儽~ꄽP   P   �섽Y넽�鄽%ꄽ�߄��愽N섽넽��섽H턽��섽�鄽+����脽�脽�脽愽�儽P   P   �焽�儽�儽�ꄽd鄽�섽j�ꄽe�Y�넽����/�l섽��m턽>턽���脽
턽P   P   �턽�鄽QꄽeꄽF턽�섽:섽s섽t鄽�섽hXꄽ�脽`섽�넽<7ꄽ>턽�脽�넽P   P   �ꄽ�鄽�넽�넽鄽w섽^愽�넽�焽�焽�넽愽儽X섽N儽<m턽�脽"鄽P   P   �섽�섽�鄽�򄽥鄽|焽��$턽������񄽌焽)섽�ℽ.焽X섽�넽��+�����P   P   X���4�焽U섽y�1儽�1.�ꄽ%�넽�ᄽ�鄽�ℽ儽`섽l섽�鄽���P   P   (넽턽V섽�ꄽ�󄽽섽��섽$넽���愽�򄽩鄽�ᄽ)섽愽�脽/��섽�P   P   �脽���������6�􄽓焽i턽���򄽺넽�焽�넽Xꄽ�����P   P   U�;턽��5��섽A����섽��]��������愽%���焽h�넽H턽~ꄽP   P   �񄽎���k�����ꄽQ턽�儽Z턽3넽������i턽���ꄽ�󄽅焽�섽Y섽OP   P   )ꄽ�愽�4턽�脽�ꄽ�ᄽ~鄽3�3넽]񄽓焽$넽.���t鄽e񄽎�8�P   P   x�ꄽ���o��섽3섽�݄��ℽ~鄽Z턽�����섽1$턽�넽s섽�ꄽ넽N턽P   P   �섽8�v��턽�ꄽ�섽&߄��݄��ᄽ�儽�섽6����^愽:섽jN섽}脽P   P   ꄽ鄽c愽�鄽v����񄽖섽3섽�ꄽQ턽A�������섽1儽|焽w섽�섽�섽�愽\턽P   P   ��넽ꄽ�����v����ꄽ�섽�脽�ꄽ�섽�󄽏�y򄽥鄽鄽F턽d鄽�߄��鄽P   P   �섽�脽�섽���鄽�턽o�4턽�5�����ꄽU섽�򄽱넽eꄽ�ꄽ%ꄽ�ꄽP   P   }脽�儽)焽�섽ꄽc愽v�����k������V섽�焽�鄽�넽Qꄽ�儽�鄽ꄽP   P   �鄽#넽�儽�脽�넽鄽8񄽖ꄽ�愽����;턽脽턽4�섽�鄽�鄽�儽Y넽焽P   P   S񄽦ㄽ�儽�䄽�߄��ㄽ�߄��܄�䄽i݄�!܄��߄�A߄�o݄��݄��ᄽ�����愽�ㄽ儽P   P   儽e䄽儽�愽�ᄽ�焽�ㄽ\܄��ℽJᄽe����䄽Zℽ�ᄽ�݄��ㄽ�愽䄽'鄽JᄽP   P   �ㄽ>ℽ�䄽u焽�䄽焽�ㄽℽㄽ�݄��߄�ބ�=ۄ��ᄽ�ᄽtᄽ$脽ZℽQᄽ'鄽P   P   �愽焽�脽�䄽Xℽ�䄽߄��ބ�iބ��ڄ����8ℽ�݄�ℽqۄ�����ބ��߄�Zℽ䄽P   P   ����|ㄽ儽�ℽ�߄��焽�ᄽp儽p愽Bㄽr䄽�儽>����愽J����߄��鄽�ބ�$脽�愽P   P   �ᄽ�ℽ����L儽�߄��儽>ᄽ�߄�.ᄽN����ᄽ�ᄽ脽�ℽ5脽ℽ�߄����tᄽ�ㄽP   P   �݄��儽�߄�]䄽ㄽ�䄽߄�wބ�4ℽ�ڄ��ℽ�ℽ�脽��䄽5脽J���qۄ��ᄽ�݄�P   P   o݄��䄽�ㄽ����܄��儽儽܄�儽����4݄�x鄽%儽焽��ℽ�愽ℽ�ᄽ�ᄽP   P   A߄�QㄽQ���Gℽ>܄�vބ��ᄽ�ބ��ᄽo��� ߄��ل��焽%儽�脽脽>����݄�=ۄ�ZℽP   P   �߄�w���ۄ��ڄ��߄��݄��݄�؄�/䄽�܄�vㄽ�ㄽ�ل�x鄽�ℽ�ᄽ�儽8ℽބ��䄽P   P   !܄�5ބ��߄��ۄ��ℽ:ڄ��ᄽ�߄��݄�Tᄽ�؄�vㄽ ߄�4݄��ℽ�ᄽr䄽����߄�e���P   P   i݄�g߄��ᄽ�܄��儽�ℽ�䄽n焽�܄�B߄�Tᄽ�܄�o��������ڄ�N���Bㄽ�ڄ��݄�JᄽP   P   䄽�ᄽw���ل��߄��䄽�鄽�儽ل��܄��݄�/䄽�ᄽ儽4ℽ.ᄽp愽iބ�ㄽ�ℽP   P   �܄�h߄��؄�݄�愽ꄽ+񄽑儽n焽�߄�؄��ބ�܄�wބ��߄�p儽�ބ�ℽ\܄�P   P   �߄�脽�߄�	ބ��ℽ�ᄽ,脽+�鄽�䄽�ᄽ�݄��ᄽ儽߄�>ᄽ�ᄽ߄��ㄽ�ㄽP   P   �ㄽI儽�ᄽ�߄��߄��؄��ᄽꄽ�䄽�ℽ:ڄ��݄�vބ��儽�䄽�儽�焽�䄽焽�焽P   P   �߄�����ᄽ�܄�/߄��߄��ℽ愽�߄��儽�ℽ�߄�>܄�܄�ㄽ�߄��߄�Xℽ�䄽�ᄽP   P   �䄽�ᄽR䄽r焽�܄��߄�	ބ�݄�ل��܄��ۄ��ڄ�Gℽ����]䄽L儽�ℽ�䄽u焽�愽P   P   �儽Qꄽ�儽R䄽�ᄽ�ᄽ�߄��؄�w����ᄽ�߄�ۄ�Q����ㄽ�߄�����儽�脽�䄽儽P   P   �ㄽm߄�Qꄽ�ᄽ���I儽脽h߄��ᄽg߄�5ބ�w���Qㄽ�䄽�儽�ℽ|ㄽ焽>ℽe䄽P   P   iՄ��؄��ل��ք��܄��ڄ��݄��܄��ބ�ۄ�܄�܄�߄��݄��߄�^ۄ�7ׄ��ք��ք�؄�P   P   ؄��ׄ��ׄ�'Ԅ�fل��ф�O݄�F߄��ׄ�$ڄ�tᄽ�ۄ��ل��ل�K݄�g܄��Ԅ�)ׄ��؄�e؄�P   P   �ք��ل�dׄ�ք�dᄽRۄ�4؄��߄��܄�`ᄽ:߄��݄�{߄�f����ڄ��ބ��؄��܄� ݄��؄�P   P   �ք��؄��ׄ��؄��؄�jք��؄�jބ�4ل��ބ�߄�Yڄ�I݄�dᄽ�܄��܄��ڄ��ׄ��܄�)ׄ�P   P   7ׄ��܄�Մ�Zۄ��ڄ��Մ�yل��ۄ��ڄ��ۄ��ڄ��ׄ��݄��ׄ�kڄ�5݄�Dۄ��ڄ��؄��Ԅ�P   P   ^ۄ������ل��ل�l߄��؄�ᄽ�݄�ل������߄�'ք��؄�?ڄ��ӄ�bℽ5݄��܄��ބ�g܄�P   P   �߄�aل�ۄ��ք��ڄ�Yڄ��؄�)ℽ-ڄ� ބ��ׄ��ڄ�vӄ�҄�vԄ��ӄ�kڄ��܄��ڄ�K݄�P   P   �݄�JՄ�>ڄ�'ᄽ�ڄ�;ބ�[ׄ��݄�S؄������ᄽ�Ԅ��܄��˄�҄�?ڄ��ׄ�dᄽf����ل�P   P   ߄�n܄�9݄��߄�jۄ�7ℽڄ�~߄��ބ��Ԅ��愽P܄��؄��܄�vӄ��؄��݄�I݄�{߄��ل�P   P   ܄�䄽�߄��ℽ7܄��ㄽ�ᄽ�ބ�e䄽�ބ�[ل�^܄�P܄��Ԅ��ڄ�'ք��ׄ�Yڄ��݄��ۄ�P   P   ܄��߄��ۄ�'܄��ބ��݄�ڄ��ڄ��܄�!ڄ�Mㄽ[ل��愽�ᄽ�ׄ��߄��ڄ�߄�:߄�tᄽP   P   ۄ�Vۄ�܄�Uℽ݄�=؄��݄�Vل�i焽�܄�!ڄ��ބ��Ԅ����� ބ������ۄ��ބ�`ᄽ$ڄ�P   P   �ބ��䄽 ބ�	䄽�����ф�>ք�Մ�h܄�i焽�܄�e䄽�ބ�S؄�-ڄ�ل��ڄ�4ل��܄��ׄ�P   P   �܄�p߄��݄��܄��؄��Є�_҄��˄�Մ�Vل��ڄ��ބ�~߄��݄�)ℽ�݄��ۄ�jބ��߄�F߄�P   P   �݄�^ӄ�Sۄ��ᄽI����ل��؄�_҄�>ք��݄�ڄ��ᄽڄ�[ׄ��؄�ᄽyل��؄�4؄�O݄�P   P   �ڄ��؄�߄�䄽܄�ᄽ�ل��Є��ф�=؄��݄��ㄽ7ℽ;ބ�Yڄ��؄��Մ�jք�Rۄ��ф�P   P   �܄��߄��܄��ބ�fׄ�܄�I����؄�����݄��ބ�7܄�jۄ��ڄ��ڄ�l߄��ڄ��؄�dᄽfل�P   P   �ք�S݄� ք�Eք��ބ�䄽�ᄽ�܄�	䄽Uℽ'܄��ℽ�߄�'ᄽ�ք��ل�Zۄ��؄�ք�'Ԅ�P   P   �ل��ք�?ׄ� ք��܄�߄�Sۄ��݄� ބ�܄��ۄ��߄�9݄�>ڄ�ۄ��ل�Մ��ׄ�dׄ��ׄ�P   P   �؄�:؄��ք�S݄��߄��؄�^ӄ�p߄��䄽Vۄ��߄�䄽n܄�JՄ�aل������܄��؄��ل��ׄ�P   P   r̄�[Ԅ��؄��Ԅ��ք�TЄ��ӄ��ք��ʄ��Є�Մ�2̈́��τ�]Ԅ��҄��Є��ք�6Մ��Ԅ��Մ�P   P   �Մ�1Մ�5؄�d҄�pք��Ԅ�Kτ��΄��ф��Є�τ��̄��҄�vф��΄�j̈́��ք��ׄ��Є�Mل�P   P   �Ԅ�Rք��ք��҄�=΄�ф��ӄ�+˄� ̈́��τ�ʄ�!τ�lτ�c˄��τ��΄�W΄��҄�/̈́��Є�P   P   6Մ�pԄ��ф�cԄ�wք�4ф�؄��҄�NՄ�aӄ��̄��Є�aф��ʄ�3ӄ��ф��Մ��ք��҄��ׄ�P   P   �ք��Є��ӄ��Є��Մ�|Ԅ�Bք��τ�r̄��̄�uτ��ӄ�|҄�cτ��ф��̈́�hɄ��Մ�W΄��ք�P   P   �Є�̈́��Մ�hՄ��τ�VЄ��̈́��̄��҄�τ�f΄�oׄ�<ф��ք�&Մ�#ф��̈́��ф��΄�j̈́�P   P   �҄�τ�QЄ��ӄ�~΄��ф�=ӄ�̈́�Zф��Ԅ�3τ�ք�eڄ�2ل�Z܄�&Մ��ф�3ӄ��τ��΄�P   P   ]Ԅ�@Մ�Є�E҄�'Մ�τ�tԄ��Ԅ��ф�ʄ��̄��τ��ӄ�߄�2ل��ք�cτ��ʄ�c˄�vф�P   P   �τ�ʄ�ф��Ȅ��΄��Ʉ��˄�̈́�̈́��Մ�˄�Sք��Є��ӄ�eڄ�<ф�|҄�aф�lτ��҄�P   P   2̈́��Ƅ�Є�τ��˄��̈́��̈́�jք�Ä�+ф�τ�dƄ�Sք��τ�ք�oׄ��ӄ��Є�!τ��̄�P   P   Մ�҄��΄�zЄ�*΄��ӄ�J̄��ф�τ��΄��ք�τ�˄��̄�3τ�f΄�uτ��̄�ʄ�τ�P   P   �Є��ф��˄�˄��˄�ф��Є�̈́�_Ȅ��τ��΄�+ф��Մ�ʄ��Ԅ�τ��̄�aӄ��τ��Є�P   P   �ʄ�dƄ��̄�7΄�Bф��܄��ل��ۄ��҄�_Ȅ�τ�Ä�̈́��ф�Zф��҄�r̄�NՄ� ̈́��ф�P   P   �ք�τ�9҄�[Є��̈́�yׄ��ڄ�SՄ��ۄ�̈́��ф�jք�̈́��Ԅ�̈́��̄��τ��҄�+˄��΄�P   P   �ӄ��҄��τ�@˄��˄�,Ԅ�N؄��ڄ��ل��Є�J̄��̈́��˄�tԄ�=ӄ��̈́�Bք�؄��ӄ�Kτ�P   P   TЄ��τ�E΄��ʄ��̈́�y҄�,Ԅ�yׄ��܄�ф��ӄ��̈́��Ʉ�τ��ф�VЄ�|Ԅ�4ф�ф��Ԅ�P   P   �ք��̈́�0ф�OЄ�Xӄ��̈́��˄��̈́�Bф��˄�*΄��˄��΄�'Մ�~΄��τ��Մ�wք�=΄�pք�P   P   �Ԅ�#Є��Մ�!Ԅ�OЄ��ʄ�@˄�[Є�7΄�˄�zЄ�τ��Ȅ�E҄��ӄ�hՄ��Є�cԄ��҄�d҄�P   P   �؄�0Є��ׄ��Մ�0ф�E΄��τ�9҄��̄��˄��΄�Є�ф�Є�QЄ��Մ��ӄ��ф��ք�5؄�P   P   [Ԅ�>ք�0Є�#Є��̈́��τ��҄�τ�dƄ��ф�҄��Ƅ�ʄ�@Մ�τ�̈́��Є�pԄ�Rք�1Մ�P   P   oӄ��ń�MÄ�Ȅ�hń��ʄ��Ä�-ń�I΄��΄��ń�_΄��΄�ń��Ä��ʄ��ń��Ȅ�QÄ��ń�P   P   �ń�>Ȅ�W�>˄��ń�9˄�B΄�Q˄��΄��Є��Ȅ�S̄��τ��ʄ�>˄��Є�1ʄ��ń��˄��ń�P   P   QÄ�/�Jń��ʄ�ʄ��Ǆ��˄��˄�Y˄�,ʄ��τ��΄�
΄��ʄ�΄�̄�vʄ�=Ƅ� ˄��˄�P   P   �Ȅ�q˄��ʄ�Ǆ�0Ȅ��Ȅ�5ń�Ą��τ�<Ǆ�X̄�L΄�˄�*̄�̄�$Ʉ�.Ǆ�uȄ�=Ƅ��ń�P   P   �ń��ń��ʄ�Ȅ�Bń�Ʉ�ʄ�	Ʉ��τ��τ�Z̄��̈́�Wń��τ��̈́��΄� ф�.Ǆ�vʄ�1ʄ�P   P   �ʄ��ʄ��Ȅ��Ʉ��Ȅ�v̈́��ʄ��̄�r̈́��Ʉ��ʄ��Ǆ�`ń��ń��Ȅ��Ä��΄�$Ʉ�̄��Є�P   P   �Ä��΄��̄��ń��ʄ�̄��ʄ��Ȅ�xτ�1Ȅ�Є��Ą����y�������Ȅ��̈́�̄�΄�>˄�P   P   ń�̈́��̈́��ń��ʄ�q΄��ʄ�Fń��̈́�Ʉ�.˄�3҄�����=Ƅ�y����ń��τ�*̄��ʄ��ʄ�P   P   �΄�@τ�:̈́��Є��ф�΄��Є�3΄�/̈́��ф��˄�Rʄ��Ȅ��������`ń�Wń�˄�
΄��τ�P   P   _΄�aЄ��˄�YȄ��Є�b˄�lɄ�˄�(ф��Ʉ��τ��҄�Rʄ�3҄��Ą��Ǆ��̈́�L΄��΄�S̄�P   P   �ń�iɄ�uф�B΄��̈́�*̄�pф��̈́�*̈́�ф������τ��˄�.˄�Є��ʄ�Z̄�X̄��τ��Ȅ�P   P   �΄��̈́��τ��΄�<΄�wȄ��Ą��҄��ʄ��ӄ�ф��Ʉ��ф�Ʉ�1Ȅ��Ʉ��τ�<Ǆ�,ʄ��Є�P   P   I΄��τ�.τ�̄�/Ƅ��Ƅ�[�����iɄ��ʄ�*̈́�(ф�/̈́��̈́�xτ�r̈́��τ��τ�Y˄��΄�P   P   -ń�˄��̄�
΄��Є��Ƅ�m����ń����҄��̈́�˄�3΄�Fń��Ȅ��̄�	Ʉ�Ą��˄�Q˄�P   P   �Ä��̄��τ�̈́�]΄��Ȅ�"���m���[����Ą�pф�lɄ��Є��ʄ��ʄ��ʄ�ʄ�5ń��˄�B΄�P   P   �ʄ��ф��̈́�ʄ��Є�#ń��Ȅ��Ƅ��Ƅ�wȄ�*̄�b˄�΄�q΄�̄�v̈́�Ʉ��Ȅ��Ǆ�9˄�P   P   hń�\Ʉ��˄�Ȅ�ӄ��Є�]΄��Є�/Ƅ�<΄��̈́��Є��ф��ʄ��ʄ��Ȅ�Bń�0Ȅ�ʄ��ń�P   P   Ȅ�Oń�YǄ�Ʉ�Ȅ�ʄ�̈́�
΄�̄��΄�B΄�YȄ��Є��ń��ń��Ʉ�Ȅ�Ǆ��ʄ�>˄�P   P   MÄ��˄��̄�YǄ��˄��̈́��τ��̄�.τ��τ�uф��˄�:̈́��̈́��̄��Ȅ��ʄ��ʄ�Jń�W�P   P   �ń�1ń��˄�Oń�\Ʉ��ф��̄�˄��τ��̈́�iɄ�aЄ�@τ�̈́��΄��ʄ��ń�q˄�/�>Ȅ�P   P   (����Ą��Ä�zĄ�qń������������t���YÄ�$������ń�������ń��Ä�Ǆ��Ä�P   P   �Ä��Ą��Ą�,Ą�����@���n���Ƅ�����¶��P�������F�������lÄ�u��������@���ń�P   P   Ǆ��Ƅ��ń�Q���Ą�zń�����)�����������ÿ��C������������Ҿ��b����ń��Ȅ�@���P   P   �Ä����Ä����ń�AÄ�4�����ξ��8���r������#���ۻ��Ժ�����1Ą��ń��P   P   ń�pń�Ӽ��8ń�cĄ�㾄�����Iń��������־��������������J�������Ą����b�������P   P   ����cĄ�п��޿���Ä�����E�����������RĄ�����\̄��Ǆ��Ä�����Ժ��Ҿ��u���P   P   �����;��ń��Ą�ܻ��&�(ń�㼄����{���Q����Ȅ��Ʉ��Ƅ��Ä�J���ۻ������lÄ�P   P   ń���������࿄�`���ƺ��j���Ä�ͼ��cƄ�MÄ�𽄽�ʄ�ń��Ʉ��Ǆ�����#���������P   P   ������������Ä�������˿��g���������������"��������ʄ��Ȅ�\̄�����������F���P   P   $���������X���񺄽X�������A���ń�Q���Ծ��.���"���𽄽Q�����������r���C�������P   P   YÄ�����B�������ҽ��H�������﹄�|��������Ä�Ծ������MÄ�{���RĄ�־��8���ÿ��P���P   P   t���y���g���8���a��ń�gĄ�𾄽�Ą�]�������Q�������cƄ�����������ξ������¶��P   P   �������O���>���u��������Ȅ�������Ą�|���ń�����ͼ��㼄��������������������P   P   ��Կ�����B���5���$ń�Ȅ��΄��𾄽﹄�A���g���Ä�(ń����Iń�4�)���Ƅ�P   P   ���м��ҽ������:����Ä��ʄ�Ȅ��Ȅ�gĄ���������˿��j���&�E�����AÄ�����n���P   P   �������Ǽ�����I���Y����Ä�$ń������ń�H���X������ƺ��ܻ������㾄�ń�zń�@���P   P   qń��Ƅ������Ä�䷄�I���:���5���u���a�ҽ��񺄽���`����Ą��Ä�cĄ����Ą�����P   P   zĄ��Ƅ������Ą��Ä��������B���>���8�������X����Ä�࿄��ń�޿��8ń��Ä�Q���,Ą�P   P   �Ä�q���������������Ǽ��ҽ�����O���g���B��������������;�п��Ӽ����ń��Ą�P   P   �Ą�BȄ�q����Ƅ��Ƅ�����м��Կ������y���������������������cĄ�pń���Ƅ��Ą�P   P   б����������1���a�������侄�C���g�������ɻ��幄�h�����������������Z�����������P   P   ����򵄽��������Z���v������� ���4����������~������A���谄�����^�������-�������P   P   ���������������粄�򷄽����	���+���b�������������»������һ��G���(���+���-���P   P   Z���x���3���#���t����Ŵ��z���ѻ��ѿ����������t���,�������Y���#���9���(�������P   P   ���N���Q���ͷ������=���򷄽۸������������������콄�N�������˸������#���G���^���P   P   ����Z�������u���G�������r�������������������&���l����������	���˸��Y���һ������P   P   ����%�������F���N���Կ��緄����������������������鰄�g�������������������谄�P   P   ���������������W�������a���V����������񷄽����I���鰄����N���,���»��A���P   P   h���򶄽Z������������������v���9�����������Ą����������l���콄�t���������P   P   幄�6��������������q���Ͼ��@���T�������C������Ą�����&��������������~���P   P   ɻ������&���Q����������R�������4Ƅ�G���kÄ�C�������񷄽�����������������������P   P   ��������[����������������������4���򺄽G���������������������������ѿ��b�������P   P   g�������������8�������ֲ��n�������4���4Ƅ�T���9������������������ѻ��+���4���P   P   C���{���k�������V���^���?������n�����������@���v���V����������۸��z���	��� ���P   P   侄����ƺ��/������;������?���ֲ������R���Ͼ������a���緄�r���򷄽Ŵ����������P   P   ��������5���񼄽�����;���^���������������q����������Կ������=����򷄽v���P   P   a�����������@�������������V���8�����������������W���N���G�������t���粄�Z���P   P   1���F������.���@���񼄽/��������������Q���������������F���u���ͷ��#�����������P   P   ����p���%����������5���ƺ��k������[���&������Z���������������Q���3����������P   P   ��������p���F��������������{���������������6���򶄽����%���Z���N���x�������򵄽P   P   o�����������&���	�������q�������C���E�������q���"������t���L�����������S��� ���P   P    ���.����������ű����������d���˱�����|�������x���������߳��ή��ί��^���\���P   P   S���X������㶄�버������������~����������E������^���*���f���z���ڱ�����^���P   P   ��������̴��<���հ���������������N���4�������騄�򫄽�������x�������ڱ��ί��P   P   ����#���쳄�֯��~���\�����������઄�����b�������ᮄ�p���2���򮄽V���x���z���ή��P   P   L���򳄽^�������>������Q�����������y���+���谄�����˶������ৄ�򮄽���f���߳��P   P   t���԰��2���ª��ڭ����������������*���Ͱ������v���_���?�������2�������*������P   P   ���V������ꪄ�����Ϭ��𫄽_�������ʦ������е��}���$���_���˶��p���򫄽^������P   P   "�������鮄������������í��5���ͯ��̳������Ĭ������}���v�������ᮄ�騄����x���P   P   q���䭄�����ݦ��������������J���a���A����������Ĭ��е������谄���������E�������P   P   ������������"���ఄ��������H���Ԭ��	�������������������Ͱ��+���b���4������|���P   P   E���.�������j������%���i���޵������3���	���A���̳��ʦ��*���y�������N����������P   P   C���ծ��c���?�����������д�������������Ԭ��a���ͯ��������������઄����~���˱��P   P   ��������㮄�����������Ӻ��鲄�����޵��H���J���5���_��������������������d���P   P   q���x�������~�������R������Ӻ��д��i�����������í��𫄽���Q�������������������P   P   ����9�������?�������R���R����������%�������������Ϭ��������\���������������P   P   	�������ִ�����������������������������ఄ�������������ڭ��>���~���հ��버�ű��P   P   &������b�����������?���~������?���j���"���ݦ������ꪄ�ª������֯��<���㶄����P   P   ����춄�寄�b���ִ����������㮄�c���������������鮄����2���^���쳄�̴���������P   P   ��������춄��������9���x�������ծ��.�������䭄�����V���԰��򳄽#�������X���.���P   P   ���������������A������֨��L������� �������G������������������S�����������/���P   P   /���w����������������������#���y���ڣ��w���X���墄�|�������v������Ť��֢��٦��P   P   ����=���Ǧ������Ħ��=���%���V�������𮄽������������߰��ᬄ���������ߩ������֢��P   P   ����������~�������m�������;������w���?���[���"���p���訄�ͤ��ת��e���ߩ��Ť��P   P   S���즄�������թ������4���j���~���ꮄ�������$���^���P�������>���ת���������P   P   ������������f���몄��������٠��D�����������"���f���c���������������ͤ������v���P   P   ��������?���:���n���N���뮄�����A��������������=���i���$�������P���訄�ᬄ�����P   P   ���u���먄�Ҩ�����^�������ū��]���q�������ש������^���i���c���^���p���߰��|���P   P   ��������9�������$���C���Ǯ��򬄽L���������������|�������=���f���$���"�������墄�P   P   G���󫄽����¬��窄�����1���⨄����[���������������ש�����"������[�������X���P   P   ����~�������$���=���7�������ë��裄����Ӭ�������������������������?�������w���P   P    ���ȭ�����뮄�`���G������ ���o����������[�������q�����������ꮄ�w���𮄽ڣ��P   P   ����V�������Y�����������p�������2���o���裄����L���]���A���D���~����������y���P   P   L���s��� �����������^�������P������� ���ë��⨄�򬄽ū������٠��j���;���V���#���P   P   ֨����������N���<�������1�������p����������1���Ǯ������뮄����4�������%�������P   P   ���4���z���f���֫����������^�������G���7�������C���^���N�����������m���=�������P   P   A���B���W���]���f���֫��<�����������`���=���窄�$������n���몄�թ������Ħ�����P   P   ������:���Y���]���f���N�������Y���뮄�$���¬������Ҩ��:���f������~�����������P   P   ����*���"���:���W���z������� ������������������9���먄�?�������������Ǧ������P   P   �������*������B���4�������s���V���ȭ��~���󫄽����u�����������즄����=���w���P   P   ���"������������������ߝ���������򞄽ݙ��(���2���R���������1�������Y���{���P   P   {���n����������M���ҡ��<���ߙ��Ĝ�������������������R���.������Ȣ�����+���P   P   Y������H������ޣ��	���O�������������疄��������������/�����������ȥ�����P   P   ��������������b���
������r���)���}������������������������y���S�������Ȣ��P   P   1�������]���_�������姄�z���{���E���̘��薄�ӛ����������|���I�������y����������P   P   ���z���؞�����
���C���ߡ��C�����������a�������󢄽_�������⥄�I������/���.���P   P   ���O���������Ɯ���������r���Q�����������ۢ��ʤ������8�������|�����������R���P   P   R�����������������p���6���P���Q���������������F���f�������_���������������P   P   2���N���F���욄�̝��V����������"���̝��@���O���J���F���ʤ��󢄽���������������P   P   (���������������������М��ݜ�����ޞ���������O�������ۢ������ӛ�������������P   P   ݙ��˗���������w���T����������!���2�����������@�����������a���薄����疄�����P   P   򞄽������������8���8�������?����������2���ޞ��̝��������������̘��}���������P   P   ����-����������d���a�����������������!������"���Q���Q�������E���)�������Ĝ��P   P   ���p���Ӛ��>���򙄽��������t�������?������ݜ�����P���r���C���{���r������ߙ��P   P   ߝ����������͞��`���ٛ��@������������������М������6�������ߡ��z������O���<���P   P   ���������������柄�f���ٛ������a���8���T�������V���p������C���姄�
���	���ҡ��P   P   ��������/����������柄�`���򙄽d���8���w������̝������Ɯ��
�������b���ޣ��M���P   P   ����z���蟄�T�����������͞��>������������������욄�����������_�������������P   P   ��������#���蟄�/�����������Ӛ����������������F���������؞��]������H�������P   P   "���3�������z���������������p���-�������˗������N������O���z�������������n���P   P   #���������������������K����������薄�q������ƙ��}���5�������З����������P   P   ����n���R���:�������đ������l���C���$���������������w������d������Ǔ��N�������P   P   ����䖄�v���e���%���J���P���b���H��������������ϛ��k���V����������.�������N���P   P   З��x�������떄�Ւ������k���A�������Л��@���̖��u���昄�����䚄�I�������.���Ǔ��P   P   ���唄�ݒ��딄�����������������������`�������瓄�V������5�������I���������P   P   �������ɔ����������h���͙������%�������@��������������5���䚄�����d���P   P   5���/���t���������������˓��򙄽h���N�������X���b����������������������V������P   P   }���	���)����G������^��������������;���2���I��������������V���昄�k���w���P   P   ƙ��[������9�������󚄽̜��&��������V���ޗ��𑄽I���b���@���瓄�u���ϛ������P   P   ���V������d���q���的�<���m����������U���Л��ޗ��2���X�����������̖����������P   P   q���u���o���䙄������������&���,���\�������U���V���;�������%���`���@����������P   P   薄�X�������m���Ӝ��<���J���(����㚄�\������������N��������Л������$���P   P   ���J�������1�������֔��(���1��� ����,��������������h��������������H���C���P   P   ��������П��/���Z���Z�������S���1���(���&���m���&������򙄽͙�����A���b���l���P   P   K���Ε��ʜ��ϔ��的������������(���J�������<���̜��^���˓��h�������k���P�������P   P   ��������A���v������-������Z���֔��<������的�󚄽������������������J���đ��P   P   ��������완�:����������的�Z�������Ӝ������q�������G���������������Ւ��%�������P   P   ��������4�������:���v���ϔ��/���1���m���䙄�d���9��������ɔ��딄�떄�e���:���P   P   �������L���4���완�A���ʜ��П����������o���������)���t������ݒ������v���R���P   P   ���򓄽����������������Ε������J���X���u���V���[���	���/������唄�x���䖄�n���P   P   <�������Ñ��+���l���鐄�����x�����������ꉄ�����F���������������&�������&���ᑄ�P   P   ᑄ�Ў������%���f�������������������v�������ˈ������􊄽���𐄽+�����Y�������P   P   &���8���Q�������挄�D���-�������a���p���=���C�������;�������-���b������-���Y���P   P   ����O���钄�o��������������O���}���k���q�������G�������G���ϊ��?���甄������P   P   &���8���䏄�����ᑄ�􎄽��������R�������ɍ������c�������i����������?���b���+���P   P   ������������"���j���0���v�������p���ꋄ�����ގ�����b���X�����������ϊ��-���𐄽P   P   ������������^�����������o�����������͌�������������Β������X���i���G����������P   P   ����މ��ڍ�����>��������������ꉄ�׍���������Д������Β��b�����������;���􊄽P   P   F���揄�������������Ԍ��ߍ������􊄽���h���F���<���Д���������c���G�����������P   P   ��������/�������(��� ���o���ކ��0���2���E���	���F����������ގ����������C���ˈ��P   P   ꉄ�����T���ꋄ�Տ�����󏄽x��������Y���E���h��������������ɍ��q���=�������P   P   ����������������z���������w���ō����������2������׍��͌��ꋄ�����k���p���v���P   P   �������u�������<�������������p���ō���0���􊄽ꉄ�����p���R���}���a�������P   P   x���֌�����獄�j�����������Ő�����w���x���ކ���������������������O�����������P   P   ����m���d���U���L���2�����������������󏄽o���ߍ������o���v�����������-�������P   P   鐄�5���=��� ���􌄽?���2����������������� ���Ԍ����������0���􎄽����D�������P   P   l���ꋄ�������K���􌄽L���j���;���z���Տ��(�������>�������j���ᑄ����挄�f���P   P   +������鐄������� ���U���獄���������ꋄ������������^���"�������o�������%���P   P   Ñ����������鐄����=���d������u�������T���/�������ڍ����������䏄�钄�Q�������P   P   ����.����������ꋄ�5���m���֌�����������������揄�މ����������8���O���8���Ў��P   