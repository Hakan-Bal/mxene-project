H   �̞�@NR>�<�`�_Rb}A?����C��8��Vb�@�w}��|A�q>��,q?Ibv�c����X��E@H            �         P   *½w½H½+½[½=½Y½�½½�½�½�½(½*½M½½�½4½E½w½P   P   w½�½�½#½;½"½>½�½�½k½�½�½^½�½}½o½)½½.½�½P   P   E½�½+½3½�½�½%½�½½½C½$½P½;½.½~½½�½�½.½P   P   4½�½�½?½/½�½�½=½�½U½�½Q½E½}½4½�½?½�½�½½P   P   �½u½�½w½Z½ ½/½7½j½½-½D½U½c½\½b½p½?½½)½P   P   ½�½i½U½�½2½W½m½ ½O½{½G½G½0½½�½b½�½~½o½P   P   M½4½X½�½T½½P½�½#½)½s½ ½�½�½�½½\½4½.½}½P   P   *½�½4½�½�½D½�½½�½:½�½B½2½�½�½0½c½}½;½�½P   P   (½½�½>½�½½�½)½½[½P½L½o½2½�½G½U½E½P½^½P   P   �½�½�½f½½-½x½d½�½�½�½½L½B½ ½G½D½Q½$½�½P   P   �½�½F½½V½e½:½½L½�½�½�½P½�½s½{½-½�½C½�½P   P   �½�½E½�½g½½½d½�½?½�½�½[½:½)½O½½U½½k½P   P   ½�½L½�½�½½�½½�½�½L½�½½�½#½ ½j½�½½�½P   P   �½L½y½½V½½>½½½d½½d½)½½�½m½7½=½�½�½P   P   Y½½�½k½P½½k½>½�½½:½x½�½�½P½W½/½�½%½>½P   P   =½½@½K½,½E½½½½½e½-½½D½½2½ ½�½�½"½P   P   [½�½U½�½�½,½P½V½�½g½V½½�½�½T½�½Z½/½�½;½P   P   +½�½f½�½�½K½k½½�½�½½f½>½�½�½U½w½?½3½#½P   P   H½�½�½f½U½@½�½y½L½E½F½�½�½4½X½i½�½�½+½�½P   P   w½�½�½�½�½½½L½�½�½�½�½½�½4½�½u½�½�½�½P   P   �½U½ ½�½�½(½�½½b½�½�½�½r½/½�½½�½�½½U½P   P   U½R½�½/½t½�½Y½�½½�½�½�½�½½�½y½�½d½0½|½P   P   ½W½½1½w½�½	½�½�½½g½�½u½'½�½�½�½�½{½0½P   P   �½�½�½�½d½�½d½�½�½�½v½�½�½q½�½�½�½[½�½d½P   P   �½Y½½O½�½�½�½�½�½�½f½`½�½^½s½�½�½�½�½�½P   P   ½�½�½�½½½o½�½�½�½�½�½�½�½�½�½�½�½�½y½P   P   �½�½�½�½�½�½�½�½�½�½�½�½�½�½�½�½s½�½�½�½P   P   /½½"½�½�½'½	½½½1½y½8½�½�½�½�½^½q½'½½P   P   r½�½�½�½Q½�½�½�½w½�½j½�½	½�½�½�½�½�½u½�½P   P   �½�½�½�½�½�½�½�½�½�½�½�½�½8½�½�½`½�½�½�½P   P   �½2½�½�½�½%½�½�½�½9½�½�½j½y½�½�½f½v½g½�½P   P   �½L½�½�½�½�½�½�½�½�½9½�½�½1½�½�½�½�½½�½P   P   b½�½�½�½P½�½ ½�½X½�½�½�½w½½�½�½�½�½�½½P   P   ½�½�½�½�½�½�½|½�½�½�½�½�½½�½�½�½�½�½�½P   P   �½	½�½�½�½�½½�½ ½�½�½�½�½	½�½o½�½d½	½Y½P   P   (½�½%½�½�½>½�½�½�½�½%½�½�½'½�½½�½�½�½�½P   P   �½�½�½�½D½�½�½�½P½�½�½�½Q½�½�½½�½d½w½t½P   P   �½Z½�½�½�½�½�½�½�½�½�½�½�½�½�½�½O½�½1½/½P   P    ½�½�½�½�½%½�½�½�½�½�½�½�½"½�½�½½�½½�½P   P   U½X½�½Z½�½�½	½�½�½L½2½�½�½½�½�½Y½�½W½R½P   P   /½M½`½C½ ½½]½J½�½½-½=½p½1½P½#½½>½k½N½P   P   N½8½�½�½�½.½w½	½$½w½�½�½l½L½½z½½�½�½�½P   P   k½½x½�½�½X½½|½½½F½v½M½�½�½r½½e½�½�½P   P   >½�½�½6½�½g½�½3½�½$½�½b½l½�½6½�½6½�½e½�½P   P   ½½½�½;½"½½*½�½:½�½�½�½�½�½4½�½6½½½P   P   #½�½�½�½�½½�½x½�½&½�½@½P½~½c½�½4½�½r½z½P   P   P½�½�½�½�½�½X½½�½5½�½a½�½=½j½c½�½6½�½½P   P   1½%½�½}½b½�½*½&½B½�½�½�½[½½=½~½�½�½�½L½P   P   p½h½P½%½�½K½A½f½�½y½G½M½½[½�½P½�½l½M½l½P   P   =½½O½½@½%½�½a½½"½w½�½M½�½a½@½�½b½v½�½P   P   -½$½½v½�½}½½�½½5½K½w½G½�½�½�½�½�½F½�½P   P   ½T½�½S½�½�½�½�½F½�½5½"½y½�½5½&½:½$½½w½P   P   �½5½�½>½0½E½½B½N½F½½½�½B½�½�½�½�½½$½P   P   J½K½2½�½�½L½f½k½B½�½�½a½f½&½½x½*½3½|½	½P   P   ]½½t½½�½�½½f½½�½½�½A½*½X½�½½�½½w½P   P   ½�½�½½*½�½�½L½E½�½}½%½K½�½�½½"½g½X½.½P   P    ½�½�½v½½*½�½�½0½�½�½@½�½b½�½�½;½�½�½�½P   P   C½½�½�½v½½½�½>½S½v½½%½}½�½�½�½6½�½�½P   P   `½�½�½�½�½�½t½2½�½�½½O½P½�½�½�½½�½x½�½P   P   M½½�½½�½�½½K½5½T½$½½h½%½�½�½½�½½8½P   P   �½�½7½�½�½v½+½]½�½�½�½�½�½4½,½�½�½�½:½�½P   P   �½�½�½�½8½�½½�½�½�½�½�½�½�½�½½�½`½�½�½P   P   :½�½C½�½F½�½�½�½½�½�½>½�½�½�½�½�½�½½�½P   P   �½�½�½�½F½�½�½�½�½�½�½�½�½�½�½�½�½�½�½`½P   P   �½<½�½.½�½�½�½�½b½�½�½�½�½�½�½�½\½�½�½�½P   P   �½�½N½g½b½{½)½�½½�½6½E½�½�½p½½�½�½�½½P   P   ,½�½�½�½�½½'½�½½�½�½f½�½	½�½p½�½�½�½�½P   P   4½�½�½�½a½�½�½@½�½�½�½�½�½�½	½�½�½�½�½�½P   P   �½�½�½�½�½�½�½�½�½�½�½�½�½�½�½�½�½�½�½�½P   P   �½½�½�½�½k½�½�½�½�½�½T½�½�½f½E½�½�½>½�½P   P   �½�½�½�½�½x½½�½�½�½�½�½�½�½�½6½�½�½�½�½P   P   �½�½#½�½½½½�½�½)½�½�½�½�½�½�½�½�½�½�½P   P   �½)½�½�½#½½t½½O½�½�½�½�½�½½½b½�½½�½P   P   ]½s½�½½½"½�½�½½�½�½�½�½@½�½�½�½�½�½�½P   P   +½�½5½�½�½½~½�½t½½½�½�½�½'½)½�½�½�½½P   P   v½½�½½q½�½½"½½½x½k½�½�½½{½�½�½�½�½P   P   �½l½�½v½�½q½�½½#½½�½�½�½a½�½b½�½F½F½8½P   P   �½6½f½�½v½½�½½�½�½�½�½�½�½�½g½.½�½�½�½P   P   7½�½�½f½�½�½5½�½�½#½�½�½�½�½�½N½�½�½C½�½P   P   �½�½�½6½l½½�½s½)½�½�½½�½�½�½�½<½�½�½�½P   P   [½½Q½½:½l½�½�½O½½�½$½?½�½�½�½½½S½½P   P   ½½½�½�½�½�½½4½�½\½1½�½K½�½�½�½�½�½½P   P   S½�½Z½�½�½½�½�½�½}½�½?½�½Q½�½�½�½½�½�½P   P   ½½½½�½½�½l½n½_½�½�½�½�½c½S½l½�½½�½P   P   ½�½M½�½3½�½�½o½k½B½½7½�½½½I½|½l½�½�½P   P   �½d½6½F½9½�½�½�½a½L½x½�½R½x½�½X½I½S½�½�½P   P   �½0½$½½5½Y½�½�½�½^½½�½�½½�½�½½c½�½�½P   P   �½4½z½U½<½_½½�½f½G½½½c½�½½x½½�½Q½K½P   P   ?½?½�½8½%½c½�½R½½�½�½�½�½c½�½R½�½�½�½�½P   P   $½I½�½J½�½�½*½�½B½X½J½:½�½½�½�½7½�½?½1½P   P   �½5½½�½�½½½�½	½*½i½J½�½½½x½½�½�½\½P   P   ½½9½`½1½'½½½T½C½*½X½�½G½^½L½B½_½}½�½P   P   O½]½½`½A½�½�½�½c½T½	½B½½f½�½a½k½n½�½4½P   P   �½&½�½�½'½½>½X½�½½�½�½R½�½�½�½o½l½�½½P   P   �½½½A½½½�½>½�½½½*½�½½�½�½�½�½�½�½P   P   l½e½p½'½�½½½½�½'½½�½c½_½Y½�½�½½½�½P   P   :½Q½½I½P½�½½'½A½1½�½�½%½<½5½9½3½�½�½�½P   P   ½r½E½�½I½'½A½�½`½`½�½J½8½U½½F½�½½�½�½P   P   Q½½N½E½½p½½�½½9½½�½�½z½$½6½M½½Z½½P   P   ½�½½r½Q½e½½&½]½½5½I½?½4½0½d½�½½�½½P   P   �½q½�½�½�½�½�½½�½�½�½�½�½"½�½�½�½�½�½p½P   P   p½b½D½�½�½�½�½#½V½½�½�½5½8½½�½�½�½�½K½P   P   �½`½½~½�½"½p½D½2½y½�½�½�½W½n½L½f½(½�½�½P   P   �½�½�½�½�½2½�½Q½�½�½�½�½n½�½�½�½Z½�½(½�½P   P   �½:½}½M½�½�½]½Y½�½�½½�½3½�½½�½½Z½f½�½P   P   �½�½�½�½�½�½�½M½�½�½½�½�½�½�½!½�½�½L½�½P   P   �½a½½�½�½�½�½½:½�½1½�½�½�½�½�½½�½n½½P   P   "½�½�½�½�½�½�½(½j½w½�½�½�½�½�½�½�½�½W½8½P   P   �½�½�½Z½|½h½�½�½x½½�½x½M½�½�½�½3½n½�½5½P   P   �½l½l½�½|½k½�½S½s½�½�½�½x½�½�½�½�½�½�½�½P   P   �½�½½�½�½�½�½½½�½z½�½�½�½1½½½�½�½�½P   P   �½�½A½�½�½�½�½�½�½Y½�½�½½w½�½�½�½�½y½½P   P   �½q½½�½�½�½½�½�½�½½s½x½j½:½�½�½�½2½V½P   P   ½�½e½�½�½�½�½�½�½�½½S½�½(½½M½Y½Q½D½#½P   P   �½�½�½�½�½�½�½�½½�½�½�½�½�½�½�½]½�½p½�½P   P   �½�½�½n½s½y½�½�½�½�½�½k½h½�½�½�½�½2½"½�½P   P   �½�½p½�½s½s½�½�½�½�½�½|½|½�½�½�½�½�½�½�½P   P   �½2½�½�½�½n½�½�½�½�½�½�½Z½�½�½�½M½�½~½�½P   P   �½�½�½�½p½�½�½e½½A½½l½�½�½½�½}½�½½D½P   P   q½d½�½2½�½�½�½�½q½�½�½l½�½�½a½�½:½�½`½b½P   P   �½.½�½½!½�½9½�½½_½�½½>½�½B½�½7½'½�½+½P   P   +½½�½�½`½�½�½�½S½l½�½½�½!½�½�½y½N½�½�½P   P   �½�½½�½�½�½½I½?½�½�½�½�½�½h½F½0½ ½�½�½P   P   '½N½,½½W½½�½�½�½4½�½p½X½½E½�½�½�½ ½N½P   P   7½½R½%½9½x½½�½½p½*½H½u½f½�½]½K½�½0½y½P   P   �½9½*½,½.½�½�½P½�½^½�½J½�½}½=½�½]½�½F½�½P   P   B½P½$½�½½b½2½�½(½'½8½H½�½[½½=½�½E½h½�½P   P   �½*½Y½�½½Z½,½�½C½�½�½I½�½g½[½}½f½½�½!½P   P   >½�½Z½A½d½7½J½ ½!½]½�½q½x½�½�½�½u½X½�½�½P   P   ½�½�½�½$½!½�½�½�½?½�½�½q½I½H½J½H½p½�½½P   P   �½�½�½�½a½2½L½�½½d½�½�½�½�½8½�½*½�½�½�½P   P   _½\½O½�½½�½�½ ½�½j½d½?½]½�½'½^½p½4½�½l½P   P   ½�½½�½½½½
½½�½½�½!½C½(½�½½�½?½S½P   P   �½½�½�½�½½�½�½
½ ½�½�½ ½�½�½P½�½�½I½�½P   P   9½I½"½�½j½�½�½�½½�½L½�½J½,½2½�½½�½½�½P   P   �½E½R½h½*½½�½½½�½2½!½7½Z½b½�½x½½�½�½P   P   !½;½*½½7½*½j½�½½½a½$½d½½½.½9½W½�½`½P   P   ½$½"½�½½h½�½�½�½�½�½�½A½�½�½,½%½½�½�½P   P   �½;½R½"½*½R½"½�½½O½�½�½Z½Y½$½*½R½,½½�½P   P   .½�½;½$½;½E½I½½�½\½�½�½�½*½P½9½½N½�½½P   P   � ½�½!½'½y½�½�½�½�½�½�½R½�½�½�½�½�½6½½�½P   P   �½�½�½�½�½½�½`½�½� ½�½½½�½m½�½½�½�½�½P   P   ½�½½�½�½½�½½�½�½½�½R½�½�½½�½,½�½�½P   P   6½w½j½/½�½&½�½6½�½�½�½�½�½�½�½�½#½x½,½�½P   P   �½r½*½�½�½½�½½|½�½½u½d½�½� ½�½�½#½�½½P   P   �½B½p½c½P½�½�½½�½�½�½�½�½{½�½�½�½�½½�½P   P   �½=½�½�½�½>½�½}½�½�½½�½�½j½�½�½� ½�½�½m½P   P   �½>½½^½z½½L½�½�½�½�½�½�½t½j½{½�½�½�½�½P   P   �½½�½w½s½d½�½	½�½� ½e½�½G½�½�½�½d½�½R½½P   P   R½�½�½�½^½]½�½�½�½^½�½�½�½�½�½�½u½�½�½½P   P   �½L½�½�½�½J½�½�½�½7½�½�½e½�½½�½½�½½�½P   P   �½A½V½�½u½5½F½s½�½X½7½^½� ½�½�½�½�½�½�½� ½P   P   �½�½�½�½u½�½�½�½�½�½�½�½�½�½�½�½|½�½�½�½P   P   �½½�½�½k½�½�½�½�½s½�½�½	½�½}½½½6½½`½P   P   �½a½b½�½�½K½�½�½�½F½�½�½�½L½�½�½�½�½�½�½P   P   �½$½ ½�½h½:½K½�½�½5½J½]½d½½>½�½½&½½½P   P   y½P½�½m½I½h½�½k½u½u½�½^½s½z½�½P½�½�½�½�½P   P   '½�½b½�½m½�½�½�½�½�½�½�½w½^½�½c½�½/½�½�½P   P   !½q½½b½�½ ½b½�½�½V½�½�½�½½�½p½*½j½½�½P   P   �½�½q½�½P½$½a½½�½A½L½�½½>½=½B½r½w½�½�½P   P   r½� ½½½� ½� ½� ½� ½� ½� ½� ½� ½� ½� ½� ½� ½� ½½� ½� ½P   P   � ½� ½ ½� ½x ½� ½� ½/½½u½� ½½n½½=½� ½� ½Z ½� ½  ½P   P   � ½� ½� ½
½!½)½� ½9½� ½x ½�½/ ½�½� ½� ½0½� ½2½ ½� ½P   P   ½� ½� ½)½Y ½½� ½½�½� ½�½� ½� ½�½� ½�½½� ½2½Z ½P   P   � ½A½� ½B½� ½� ½� ½½½� ½l½Z½M½f½p½� ½� ½½� ½� ½P   P   � ½� ½� ½� ½� ½� ½� ½4½�½� ½½½2½½½½� ½�½0½� ½P   P   � ½5½� ½� ½� ½)½� ½C½� ½� ½k½½2½�½M½½p½� ½� ½=½P   P   � ½� ½%½� ½� ½½� ½� ½� ½� ½�½h½.½�½�½½f½�½� ½½P   P   � ½p ½� ½
½� ½� ½½R ½� ½�½�½� ½4½.½2½2½M½� ½�½n½P   P   � ½� ½� ½� ½� ½� ½� ½� ½� ½� ½ ½. ½� ½h½½½Z½� ½/ ½½P   P   � ½½� ½� ½� ½½� ½� ½½"½
½ ½�½�½k½½l½�½�½� ½P   P   � ½'½� ½� ½� ½5½#½� ½� ½� ½"½� ½�½� ½� ½� ½� ½� ½x ½u½P   P   � ½� ½� ½� ½� ½� ½� ½� ½� ½� ½½� ½� ½� ½� ½�½½�½� ½½P   P   � ½Z ½� ½� ½� ½� ½] ½t ½� ½� ½� ½� ½R ½� ½C½4½½½9½/½P   P   � ½� ½� ½� ½� ½!½� ½] ½� ½#½� ½� ½½� ½� ½� ½� ½� ½� ½� ½P   P   � ½5½#½½� ½½!½� ½� ½5½½� ½� ½½)½� ½� ½½)½� ½P   P   � ½� ½� ½� ½� ½� ½� ½� ½� ½� ½� ½� ½� ½� ½� ½� ½� ½Y ½!½x ½P   P   ½Q½� ½� ½� ½½� ½� ½� ½� ½� ½� ½
½� ½� ½� ½B½)½
½� ½P   P   ½� ½� ½� ½� ½#½� ½� ½� ½� ½� ½� ½� ½%½� ½� ½� ½� ½� ½ ½P   P   � ½� ½� ½Q½� ½5½� ½Z ½� ½'½½� ½p ½� ½5½� ½A½� ½� ½� ½P   P   ���� ½� ½? ½� ½� ½����L ½~ ½@ ½! ½ ½b ½# ½����� ½{ ½@ ½� ½ ½P   P    ½' ½� ½����( ½. ½: ½t ½� ½� ½; ½ ½t ½� ½� ½2 ½N ½' ½����� ½P   P   � ½����� ½ ½# ½f ½. ½B ½c ½� ½k ½½� ½� ½? ½H ½ ½] ½  ½����P   P   @ ½��������H ½ ½V ½X ½� ½ ½� ½����� ½� ½����� ½- ½� ½j ½] ½' ½P   P   { ½����q ½����o ½e ½ ½� ½ ½f ½� ½
 ½½����� ½� ½����� ½ ½N ½P   P   � ½D ½u ½a ½Z ½� ½ ½W ½����u ½� ½n ½� ½� ½r ½w ½� ½- ½H ½2 ½P   P   ����R ½����. ½ ½; ½ ½z ½n ½� ½� ½e ½� ½. ½� ½r ½� ½� ½? ½� ½P   P   # ½| ½! ½U ½[ ½ ½w ½0 ½� ½� ½���� ½� ½( ½. ½� ½��������� ½� ½P   P   b ½� ½ ½ ½J ½ ½A ½� ½� ½� ½g ½� ½½� ½� ½� ½½� ½� ½t ½P   P    ½x ½. ½H ½V ½h ½0 ½M ½z ½1 ½& ½½� ½ ½e ½n ½
 ½� ½½ ½P   P   ! ½f ½- ½P ½����2 ½  ½( ½+ ½� ½4 ½& ½g ½����� ½� ½� ½����k ½; ½P   P   @ ½� ½� ½I ½M ½0 ½ ½} ½` ½_ ½� ½1 ½� ½� ½� ½u ½f ½� ½� ½� ½P   P   ~ ½� ½ ½> ½� ½x ½����g ½h ½` ½+ ½z ½� ½� ½n ½���� ½ ½c ½� ½P   P   L ½� ½I ½; ½~ ½> ½� ½� ½g ½} ½( ½M ½� ½0 ½z ½W ½� ½� ½B ½t ½P   P   ����` ½B ½/ ½ ½  ½# ½� ½���� ½  ½0 ½A ½w ½ ½ ½ ½X ½. ½: ½P   P   � ½f ½) ½ ½V ½D ½  ½> ½x ½0 ½2 ½h ½ ½ ½; ½� ½e ½V ½f ½. ½P   P   � ½R ½����N ½_ ½V ½ ½~ ½� ½M ½����V ½J ½[ ½ ½Z ½o ½ ½# ½( ½P   P   ? ½����h ½T ½N ½ ½/ ½; ½> ½I ½O ½H ½ ½U ½. ½a ½����H ½ ½����P   P   � ½����� ½h ½����) ½B ½I ½ ½� ½- ½. ½ ½! ½����u ½q ½����� ½� ½P   P    ½������������R ½f ½` ½� ½� ½� ½f ½x ½� ½| ½R ½D ½������������' ½P   P   ����s���L���O�������r�������������������5 ½ ½��������������������G���Q���t���P   P   t���}���_���e�������a���9 ½����O���*��� ½��������o�������  ½���� ½\���i���P   P   Q�������M���f�������u���������������c ½y���! ½����z ½������������\�������\���P   P   G�����������E��� ½b���x�����������- ½ ½������������# ½������������\��� ½P   P   �����������
�������������������t ½ ½����W ½����B ½ ½, ½H ½������������P   P   ��������z���z�������~��� ½����o���) ½����6 ½ ½ ½Q ½B���, ½��������  ½P   P   ����W���������������9���������������L ½����> ½� ½I ½g ½Q ½ ½# ½��������P   P   ��������v�����������������������Q���S ½ ½^ ½ ½+ ½I ½ ½B ½����z ½o���P   P   ��������R����������x���O�����������,��������������� ½� ½ ½����������������P   P    ½����s������������������������������� ½1 ½����^ ½> ½6 ½W ½����! ½����P   P   5 ½���������������`���x�������i���0���P ½ ½���� ½������������ ½y��� ½P   P   ����9�������f���e�����������������������0�������,���S ½L ½) ½ ½- ½c ½*���P   P   ��������j���h������[���R���O�����������i�����������Q�������o���t ½��������O���P   P   �����������������������(���A���O�����������������������������������������������P   P   ��������e�������|�����������(���R�������x�������O����������� ½����x�������9 ½P   P   r���[�������y�������y����������[�������`�������x�������9���~�������b���u���a���P   P   ����������������&�������|����������e������������������������������ ½��������P   P   O�������m�����������y�����������h���f�����������������������z���
���E���f���e���P   P   L�����������m�����������e�������j�����������s���R���v�������z�����������M���_���P   P   s�������������������[���������������9������������������W������������������}���P   P   ��������g��������������5���,���L���@�������_���O���'���1���������������h�������P   P   �������������������}�����������S�����������������S������������������� �������P   P   h�������i�������������Y������3���$���������������7������)���\����������� ���P   P   �����������������������K�����������c�������L���S�������l�����������d�����������P   P   ����+���^���#�����������X�������?������H�������/�������<���5���G�������\�������P   P   ����K�����������[�����������$���l���K�������?���^���Z���Y�������5�������)�������P   P   1����������R�����������)�������-����������N���������������Y���<���l����������P   P   '�������!�����������K������&���Q���������� ½a�����������Z�����������7���S���P   P   O����������2��������������r���T�����������T������a�������^���/���S�����������P   P   _�����������������������������������;���
�������T��� ½N���?�������L����������P   P   �������V���������������q�������+���#�������
������������������H��������������P   P   @���3���Z������������������� �������`���#���;��������������K������c���$�������P   P   L�������5�������F�������������������+�������T���Q���-���l���?�������3���S���P   P   ,���~������������������������������ �����������r���&�������$������������������P   P   5��������������u���������������������q��������������)�������X���K���Y�������P   P   ��������5����������������������������������������K����������������������}���P   P   ����V�������������������u�������F���������������������������[�������������������P   P   ����������Q����������������������������������2�������R�������#������������P   P   g�������������������5�����������5���Z���V����������!�����������^�������i�������P   P   ���������������V����������~�������3���������������������K���+���������������P   P   '�����������&�����������T���<���C���)���Q������F���f���H��������������������P   P   ����������*�����������a���a�������U�����������g�������Z���d�����������������P   P   ���$��������������v������Z��������������&�������*�������b������^���������P   P   �����������1������h����������#���4�������������������9������}���7���^�������P   P   �����������������������"������������������D���V���^�������������}����������P   P   ��������N���N�����������k���P����������������������\������������������b���d���P   P   H���	�������������������3���a�������B����������B������o����������9�������Z���P   P   f����������!���1������� ���c������� �������q���|���+������\���^�������*�������P   P   F���j���s�������^�������V���y���0���X��������������|���B�������V�����������g���P   P   ���S���������������������������V���'��������������q�����������D�������&�������P   P   Q���w�������,�������I���c���?�������j���D�������������������������������������P   P   )���n�����������/���z�������"�����������j���'���X��� ���B�����������4������U���P   P   C���B����������@��������������G�����������V���0������������������#�����������P   P   <�����������<����������&�����������"���?�������y���c���a���P�����������Z���a���P   P   T���*���U�������l�����������&����������c�������V��� ���3���k���"���������a���P   P   ��������������������0���������������z���I���������������������������h���v�������P   P   ������������3���H�������l������@���/�����������^���1��������������������������P   P   &�������L�������3�����������<�����������,�����������!�������N�������1������*���P   P   ������������L�����������U����������������������s�����������N������������������P   P   ����;�������������������*�������B���n���w���S���j������	���������������$������P   P   x���=�������U������a���S���k�������"���1���������������=���C���7���P���.���@���P   P   @���F�������?���[���H�������!�������������8���������� �������G���C���)�������P   P   .���*�������������j���b�������i���)���������������6�����������J���d�������)���P   P   P���W���q���\���h���w�����������D�����������7���9�������}���?�����������d���C���P   P   7���u�������l������2���Y�������\���"���<���I�������p���N������y�������J���G���P   P   C���6���������R���[�����������X��������������Y���'���n����������?�����������P   P   =����������������������B������v���q���i���}����������3���n���N���}������� ���P   P   ������������/���=�������������������N�������Z���D���Q������'���p�������6�������P   P   ��������^��������������k�������������������N�������D�������Y�������9����������P   P   �����������\���������]��������������8�������N���Z���}�������I���7�������8���P   P   1�������T���3���x���
���~���V���i����������8�����������i�������<��������������P   P   "������������������d���q��������������������������N���q������"�������)�������P   P   ��������{�����������W�������j���!�������i���������������v���X���\���D���i������P   P   k�������
���4�������������������j�������V����������������������������������!���P   P   S�������J���V�������~���������������q���~���]���k�������B�������Y�������b�������P   P   a���������������)�������~�������W���d���
������������������[���2���w���j���H���P   P   ���D�������L���K���)������������������x���������=�������R������h�������[���P   P   U���|���#������L�������V���4�����������3���\�������/���������l���\������?���P   P   ����o�������#�����������J���
���{�������T������^������������������q����������P   P   =���F���o���|���D�������������������������������������������6���u���W���*���F���P   P   O������l���R������������������������������������$�������~�������N����������P   P   ���������������������������>���+����������%����������&����������������������P   P   �����������{���<�������L�������g�������������������������������8�������?�������P   P   N�����������B�����������������3���d���}�����������o���W���5������������������P   P   ����o���<���b����������B����������������������������������d�����������8�������P   P   ~�������8���4�������k�����������]���U�������������������j������d���5����������P   P   ����q���x�����������w�������+���j���B�������|�����������$���j�������W�������&���P   P   $�������8���2���$���#�����������������m���{����������������������o����������P   P   �������i�������T������������������v�����������������������������������������P   P   �������������������t�����������������)�����������{���|�������������������%���P   P   ����������������/���W���I������� �����������)�������m���������������}����������P   P   �������x���q���Q���#���!���(���]��������������v�������B���U�������d�����������P   P   ����������u���K���������������w���]��� ������������j���]�������3���g���+���P   P   ������������~���3�������&���$�������(������������������+�������������������>���P   P   ��������_�������R���$�������&�������!���I�����������������������B������L�������P   P   ����o���)�����������A���$�����������#���W���t�������#���w���k������������������P   P   ������������=���1�������R���3���K���Q���/�������T���$������������������<�������P   P   R���w���P���`���=�����������~���u���q���������������2�������4���b���B���{�������P   P   l����������P�������)���_����������x�����������i���8���x���8���<���������������P   P   ����������w�������o����������������������������������q�������o��������������P   P   ����)�������?�������+�������e���R�������3�������\���[�������.���v���9�������(���P   P   (���������\�������
�����������`�������������������b�������������������k�������P   P   ������������_��������������i���"��������������,�������&���R���/�������a���k���P   P   9�����������$�������������������d���X���E���|���q���N���\���n�������m�����������P   P   v���Y�������O�����������.���������������b�������,�������b���������������/�������P   P   .���s�����������F����������H�������������������=���c���������������n���R�������P   P   ������������.�������������������$���M���p����������	�����������b���\���&�������P   P   [������������������������L���r�������V�������?������	���c�������N�������b���P   P   \�����������p���f���������������_�������5���_���^���?������=���,���q���,�������P   P   �����������g�������f���N����������������������_�������������������|�����������P   P   3���������������d�������x���������������?�������5���V���p�������b���E����������P   P   ��������������������������������������������������������M�����������X�����������P   P   R������������������� ���������������������������_���r���$�����������d���"���`���P   P   e������������������������������������������������L�������H�����������i�������P   P   ����
�������l���`�����������������������x���N������������������.��������������P   P   +���������������h������������� �����������f������������������������������
���P   P   ����F�����������x���h���`���������������d�������f�����������F�������������������P   P   ?���h�������	�����������l�������������������g���p������.�������O���$���_���\���P   P   ������������������������������������������������������������������������������P   P   )�����������h���F�������
����������������������������������s���Y��������������P   P   l���;���G����������������������)�������]����������U���-�������g����������:���P   P   :���'���A���d����������������h���e���O���&���Y�������#�����������.�������L���P   P   �������:���{���m�������t�����������i���������������I��������������������������P   P   ����"����������	�����������n���2�����������{���������������C���n���q�������.���P   P   g��������������������������Z���������������?���m������������������n�����������P   P   �������G���j�������������������E������������������O���������������C�����������P   P   -�������������������������������������������w�������"�������������������#���P   P   U�������A���J���'���-�������k�������%���������������������O����������I�������P   P   ���%�������`���������������!������`�������[����������v������m�����������Y���P   P   ����[�������������������������L������� ��� ���[��������������?���{�������&���P   P   ]��������������9�������O�����������#���V��� �������������������������������O���P   P   ����=�����������Z���a���b���P�����������#�������`���%�������������������i���e���P   P   )���������������V���J�������=���g�����������L�������������E�������2�������h���P   P   ����������������l���A�����������=���P����������!���k����������Z���n����������P   P   �����������������Q���������������b���O������������������������������t�������P   P   �������3���Q�����������Q���A���J���a���������������-�������������������������P   P   ������������8��������������l���V���Z���9�����������'���������������	���m������P   P   ��������^�������8���Q���������������������������`���J�������j�����������{���d���P   P   G���������^�������3�����������������������������A�������G���������:���A���P   P   ;���������������������������������=������[���%������������������"�������'���P   P   ������Z���`��������������������������=���*���k�������$�����������c���1�������P   P   �������������������A�������I�����������������������;���J�������@��������������P   P   1���G���H�������Z���P�������e������;�������C��������������g�������a���?������P   P   c���~���W���m�������T��������������g���m���>���I�������q����������}���a�������P   P   ����m���������������C�����������N����������R�����������������&�����������@���P   P   ����������������������������g��������������R���:���{���{��������������g�������P   P   $�����������D���������������9������j���	���n����������i���{������q�������J���P   P   ������������������������z�������0�������������S����������{�������������;���P   P   k�����������B�������]�����������O�����������$���0���S�������:�������I�����������P   P   *������������������d���������������C�������k���$������n���R���R���>���C�������P   P   =������������������,�����������	����������������������	����������m�����������P   P   ����������������������������|�����������C����������j�����������g���;�������P   P   ����/�������v���R���x���$���n���k���|���	�������O���0���������N�������������P   P   ����������������+���w�����������n����������������������9���g�����������e���I���P   P   ���o�������������������:�������$������������������z���������������������������P   P   ���������������q���`�������w���x������,���d���]���������������C���T���P���A���P   P   �������������������q�������+���R��������������������������������������Z�������P   P   `���e�������`������������������v���������������B�������D�����������m�����������P   P   Z���l������������������������������������������������������������W���H�������P   P   ���0���l���e�����������o�������/������������������������������m���~���G������P   P   ��������9��������������������������������������|���g������������������4���{���P   P   {������a�����������	���c����������U����������b�����������a��������������p���P   P   4�������B�����������8����������}���t���E���Z���V���M���������������C�����������P   P   �����������������Y�������8�������b�������������������m�������F������C�������P   P   ��������(������������������9�������)�������W�������8�������0�������F����������P   P   ����=������ ���1�������W�����������������&���!���D���<������0�����������a���P   P   ������������������������������[���]�������5���=����������<�������m�����������P   P   g���u����������3���}���S���x�������t�������(���0�����������D���8�������M�������P   P   |���_����������������������r���]���W��� ����������0���=���!�����������V���b���P   P   ������������O�����������K���������������������������(���5���&���W�������Z�������P   P   �����������������������������$�������������� ����������������������E������P   P   ���������������������������������������������W���t���]������)���b���t���U���P   P   ���������������,���~���"���~���:�������$�������]�������[���������������}�������P   P   ����P�������������������
������~���������������r���x�����������9���8����������P   P   ����W���
���M�����������$���
���"�����������K�������S�������W��������������c���P   P   �������������������u�����������~������������������}�������������Y���8���	���P   P   ����R�������%���7���������������,�����������������3�������1�������������������P   P   ����������<���%�������M�������������������O������������� ������������������P   P   9�������?��������������
������������������������������������(�������B���a���P   P   ����������������R������W���P�����������������_���u�������=�����������������P   P   �������O�������"�����������+���"���l���|���/���<���:���|�������?�������J�������P   P   ��������+�������A���5���m������r����������������P������r���$���%�������7���P   P   J���.���\�����������$������}�����������n���m���e��������������� ���*����������P   P   ��������������-���@�������[���Q���A�����������������Q���)���E�������*���%���P   P   ?��������������9���(������<������� �������������������z����������E��� ���$���P   P   ����Q����������M�������]�������X���/���	���7���1���#���6���������)�������r���P   P   |����������������������������������8������8���������������6���z���Q����������P   P   :���B�������������������0���!���a��������������.�����������#��������������P���P   P   <���H�������J��� ���%�������_���*�������D�����������.�������1�����������e������P   P   /�����������1���%���@���D���\�������E������u�����������8���7�����������m������P   P   |�������6���'���H�������,���)���N�������n������D���������	����������n������P   P   l�����������������{���~������������������E�����������8���/��� ���A�����������P   P   "�������W������W���U���
���^���G������N�������*���a�������X�������Q�������r���P   P   +���k��������������l�����������^�������)���\���_���!����������<���[���}������P   P   ����F�������/���s���������������
���~���,���D�������0�������]�������������m���P   P   ������������U���=���L�������l���U���{�������@���%���������������(���@���$���5���P   P   "���`���������������=���s�������W�������H���%��� �����������M���9���-�������A���P   P   �������������������U���/������������'���1���J������������������������������P   P   O������������������������������W������6�����������������������������\���+���P   P   ���2���������`�������F���k�������������������H���B�������Q����������.�������P   P   B���������������������������c���������������{���������������{�������������������P   P   ��������T�����������l������L���$�������B���������������<�������M�����������a���P   P   ����/������������������@�������\������D���I���������~�������c��������������P   P   ����v���u�������������������W�������*���"���D���4���.���.�������0���������������P   P   ����!�������*�������Y���h���.�������5�������&�������U�������-�������0���c���M���P   P   {���a�����������j���y���������������T������� ½ ½G ½��������-���������������P   P   ����q���\���1���]���[�������S���^����������  ½� ½q ½� ½��������.���~���<���P   P   ����������������������������`�������4������]���o ½� ½q ½G ½U���.����������P   P   ��������R��������������D���������������/���V���e���o ½� ½ ½����4����������P   P   {�����������K���"���C���i���k�������{���n������V���]���  ½ ½&���D���I�������P   P   ����7�������W����������\���W��������������n���/������������������"���D���B���P   P   �������e�������O���!���2���\�������s������{�������4������T���5���*����������P   P   ��������������������N�������T���������������������������^���������������\���$���P   P   c����������F���9���]�����������T���\���W���k�������`���S�������.���W�������L���P   P   �����������N�������F���b�����������2���\���i���D���������������h�������@������P   P   ����c�����������A�������F���]���N���!������C�����������[���y���Y�����������l���P   P   ����m���m�����������A�������9�������O�������"����������]���j������������������P   P   ����U�������C�����������N���F�����������W���K�����������1�������*���������������P   P   ����w�����������m������������������e�����������R�������\�����������u�������T���P   P   �������w���U���m���c�����������������7���������������q���a���!���v���/�������P   P   ���������������A�������j���n�������'�������������������w�������?���������������P   P   ������������-���1�������&�����������s�����������s���u��������������"���@�������P   P   ����s�������Q�������D�������k������� �����������c���=�������f�������4�������@���P   P   ����|�����������#���!�������N���������������]���U�������p�������J�������4���"���P   P   ?���������������+�����������U��������������� ½M½
½�����������J�����������P   P   ����F�����������i����������V�������'���M ½�½�½�½~½u ½�������f������P   P   w�������I���t���8�������q����������q��������½T½Q½�½~½����p�����������P   P   ��������,�����������9�������r���_���+�������½�½v½Q½�½
½����=���u���P   P   ����2�������Z�������O��������������m�������s���½�½T½�½M½U���c���s���P   P   ������������7�����������B�������������������k���s���½�½�½� ½]�����������P   P   ����z���z�������W�������H�������a���e�����������������������M ½����������������P   P   '���w������.�������<���A�������*������e�������m���+���q���'���������� ���s���P   P   ����[�������:���N�������W�������>���*���a�����������_��������������������������P   P   n���P���������������������������������������������r�������V���U���N���k�������P   P   j�����������6���c���L���X�������W���A���H���B�����������q������������������&���P   P   ��������,��������������L�����������<�����������O���9���������������!���D�������P   P   A���`���I�������W������c�������N�������W���������������8���i���+���#�������1���P   P   ������������������������6�������:���.�������7���Z�������t���������������Q���-���P   P   ���������������I���,�����������������z�����������,���I�����������������������P   P   ����h�����������`�����������P���[���w���z�������2�����������F�������|���s�������P   P    ������n����������S���l���'���&���������������������h���Y������������������P   P   �������j���7���L��������������2������������������=�����������,���J���,���X���P   P   �������S���8�������������������������������������C���d�������m����������,���P   P   ����������������P����������I�������1���� ½d½`½� ½������m���*�������J���P   P   ����N�������0�������<���g�������2�������½ ½�½4½½ ½����m���m���,���P   P   Y�������������������[�������������������9½½�½�½½*½ ½�����������P   P   h���1����������������c�����������8���½½�½g½�½½½���d�������P   P   ������p�����������m������"���������r ½%½�½r½g½�½4½� ½C���=���P   P   ���������������������������R���6����������g½�½�½�½�½�½`½��������P   P   �����������q���e���S���Z������������������_���g½%½½½ ½d½��������P   P   ������������Y��������������4�����������������������r ½½9½½� ½��������P   P   ��������X���������������������������B�����������������8�����������1���������P   P   &����������������������������������������������6��������������2�����������2���P   P   '�����������M��������������������������4�������R���"���������������I�����������P   P   l����������h�����������
������������������Z����������c�������g��������������P   P   S���F���o�������p���������������������������S�������m������[���<��������������P   P   ������������������p����������������������e�����������������������P������L���P   P   �����������(�����������h���M�����������Y���q������������������0�������8���7���P   P   n�����������������o���������������X���������������p������������������S���j���P   P   ���1��������������F��������������������������������1�������N��������������P   P   .���,�����������M�����������'�������3�������z�����������b������������������*���P   P   *���=��������������J���O�������_�������
�������I�����������-���j�������i�������P   P   ����5�������n�������������<�����������w ½� ½� ½��������9���������������i���P   P   �������� ���������������j����������� ½�½�½�½h½� ½;�������������������P   P   ���>�������&������o���������������½8½�½�½�½E½�½������������j���P   P   ����*�����������?�������)���Q��������½�½�½�	½�	½�½�½�½;���9���-���P   P   b���������J����������h�����������)½½�½�
½�
½�
½�½E½� ½��������P   P   �������������������������������L�������t½�½�	½b
½�
½�	½�½h½��������P   P   ����������������������������@�������q���v ½�½�½�	½�
½�	½�½�½� ½I���P   P   z���w���V������M���N�������{���h���%�������� ½�½�½�½�½�½�½� ½����P   P   ����������������|�������������������#�����������v ½t½½�½8½�½w ½
���P   P   3���E���9���Y�������?����������_�������#���%���q�������)½�½�½� ½��������P   P   ������������I�������5����������P���_�������h�������L���������������������_���P   P   '���i���|���������������m������������������{���@����������Q�����������<�������P   P   ��������������������������m��������������������������h���)�������j������O���P   P   ���������������Z�������������5���?�������N�������������������o����������J���P   P   M���E���,�����������Z�������������������|���M��������������?������������������P   P   �����������N������������������I���Y������������������J�������&�������n�������P   P   ���������������,�����������|�������9�������V���������������������� ����������P   P   ,���j���������E����������i�������E�������w��������������*���>�������5���=���P   P   W���������������`�������������������p��������������U�����������B���f�����������P   P   ������������5���t�����������q�����������z���E���z�����������������������������P   P   �������������������������u�������7½�½�½�½L½@���q�����������������P   P   f���������f���������������a��������½5½?	½Z	½½�½����K��������������P   P   B�������2�������P�����������h���e ½½
½g½E½Q½.
½3½S ½K�����������P   P   ����.���l���e���.�����������u�������K½½{½�½�½�½�
½3½����q�������P   P   ����)���w������������������n���f����½�	½�½/½�½½�½.
½�½@�������P   P   U���Y�������?���.�������S���U���}���½"½�½�½h½�½�½Q½½L½����P   P   �������H���u�������^���D���������������|½:	½½�½/½�½E½Z	½�½z���P   P   ����k���V���G�����������:���c���_���k���D����½:	½�½�½{½g½?	½�½E���P   P   ���&���������������#���y���`�������C������D���|½"½�	½½
½5½�½z���P   P   p���i���������������g���U�����������n���C���k�������½�½K½½�½7½����P   P   ��������������������o������`���?�����������_�������}���f�������e ½������������P   P   ���� ���c�����������E�����������`�������`���c�������U���n���u���h���a���u���q���P   P   ����`�������b�������e���@����������U���y���:���D���S���������������������������P   P   ����"������`�������]���e���E���o���g���#�������^������������������������������P   P   `���B�������F���9�����������������������������������.�������.���P����������t���P   P   ��������~�������F���`���b�������������������G���u���?�������e�������f������5���P   P   �������K���~��������������c���������������V���H�������w���l���2��������������P   P   ����E����������B���"���`��� �������i���&���k������Y���)���.�����������������P   P   ��������^���h�����������������������������������������������������U���<�������P   P   ������������Z���B���\������j���"��������½y½�������E������:���$���J�������P   P   <�������Y���Q�������+����������� ½l½l½�½i½n½� ½��������������J���P   P   U����������O���A������r���`����½v	½\½�½�½>½\	½t½8����������$���P   P   �������d����������)�������F����½½2½1½9½%½X½½�½8�������:���P   P   ����h�����������l��������������x½*½�½�½'½½�½�½½t½������P   P   ����t����������r���T�������C���� ½b	½½~½½�½/½�½X½\	½� ½E���P   P   ��������������������������������
���C½H½?½ ½�½�½½%½>½n½���P   P   ����m�������V��� ���$�������o�����������V½�½
½ ½½'½9½�½i½����P   P   ��������d�������������������M���z���t���p½�½�½?½~½�½1½�½�½y½P   P   �������W����������J�������	���*�����������p½V½H½½�½2½\½l½�½P   P   �����������q���Y���S���_���`���f�����������t�������C½b	½*½½v	½l½����P   P   ��������N���u���[������������������f���*���z�������
���� ½x½�½�½� ½"���P   P   ����y���W���?���`�������R���&�������`���	���M���o�������C�������F���`������j���P   P   �����������������������y���R�������_������������������������������r����������P   P   ����x�������7�������a���������������S���J�������$�������T�������)������+���\���P   P   ����������������V�����������`���[���Y����������� �������r���l�������A�������B���P   P   h���B�������	�������7�������?���u���q����������V������������������O���Q���Z���P   P   ^������u������������������W���N�������W���d������������������d�������Y�������P   P   �����������B�������x�������y�������������������m�������t���h�����������������P   P   n���L������������������T����������R�������,���������5�����������s�������@���P   P   @���F���
���B��������������r�������½�½�½�½��������������Z���/���
���P   P   ������������;�����������>��� ���+½�
½�½�½�½o
½e½��������������/���P   P   s�����������y�����������D���(����½�½½�½�½ ½½�½���C�������Z���P   P   ����+�������;�����������2������b	½0½F½&½�½.½r½
½�	½����������P   P   ���������������������������������½�½c½5"½�$½�$½"½x½
½�½������P   P   5���H�������v�������,���0���3���+½]½�½"½h&½)½�&½"½r½½e½���P   P   ����������!���4���;���������������v
½�½½�$½7)½)½�$½.½ ½o
½����P   P   ������������������������������������½�½u½ ½�$½h&½�$½�½�½�½�½P   P   ,����������������������.�����������7���y½�½u½½"½5"½&½�½�½�½P   P   ������������i�������$�������z�������`���f���y½�½�½�½c½F½½�½�½P   P   R���z���:���P������������������(���0���`���7����½v
½]½�½0½�½�
½�½P   P   �����������_����������������������(�������������������+½�½b	½�½+½���P   P   ���0���������������)�������������������z���������������3����������(��� ���r���P   P   T���)���
���W�������C���������������������.�����������0�������2���D���>�������P   P   ����^���_�������������C���)�����������$�����������;���,����������������������P   P   �����������`��������������������������������������4���������������������������P   P   ����n�����������`�������W�������_���P���i����������!���v�������;���y���;���B���P   P   �������������������_���
����������:��������������������������������������
���P   P   L�����������n������^���)���0�������z�������������������H�������+�����������F���P   P   u���a�������x���h���B���=�����������f�������������������������Y���]�������R���P   P   R���Z�����������D����������I����½_½�½�½[½s½���*���h���������������P   P   ����@�����������v�������9���k���W
½�½�½8½�½�½{
½>����������q�������P   P   ]�����������n����������i����½�½?½� ½�$½�$½� ½3½�½y½K�����������P   P   Y���������������J���i������k½½�½�&½%-½c/½1-½�&½�½½y½���h���P   P   ����+�������~���1���������:���
½�½�(½?1½D6½T6½1½*)½�½�½>���*���P   P   �����������<������������������&
½�½9'½+1½�7½R;½�7½1½�&½3½{
½���P   P   ����m�������q���x�������V��������½�½� ½�,½.6½w;½R;½T6½1-½� ½�½s½P   P   ����K������S���Q���H������i���j���½}½�$½�/½.6½�7½D6½c/½�$½�½[½P   P   �����������������
���������������9���m½%½�$½�,½+1½?1½%-½�$½8½�½P   P   ����h���������������D����������������������m½}½� ½9'½�(½�&½� ½�½�½P   P   f���4�����������9���0���F�������j����������9���½�½�½�½�½?½�½_½P   P   ����������������M���"������(���j���j�����������j����½&
½
½½�½W
½�½P   P   ������������������s����������(���������������i����������:���k½�½k���I���P   P   =������������������y�������������F��������������V�������������i���9������P   P   B���������������_���L���y���s���"���0���D���
���H��������������i���������������P   P   h���]�����������X���_����������M���9����������Q���x�������1���J������v���D���P   P   x���8�������b�����������������������������������S���q���<���~�������n�����������P   P   ����������������������������������������������������������������������������P   P   a���V�������8���]�������������������4���h�������K���m�������+�����������@���Z���P   P   ����b���������������������������
���y ½½9 ½����{���6�������`�����������O���P   P   O���F���2���i�������c���h���h����½�½
½ ½�½�½C���E���
�������J�������P   P   ����N�������V�������Z���'����½?½�½�#½/&½�#½�½#½Y½���Q���o���J���P   P   ����w���������������h�������½�½�%½�0½�5½y5½�0½�%½�½�½����Q�������P   P   `��������������������������½Q½�*½A8½@A½�C½:A½�7½�*½_½�½���
���P   P   ��������w���|�������w���U���Z½�½�*½�:½tG½�M½N½�G½�:½�*½�½Y½E���P   P   6���N����������$���l���"���<����½�%½48½�G½ZQ½	S½;Q½�G½�7½�%½#½C���P   P   {���	�������!������R�������W����½�½�0½	A½�M½�R½	S½N½:A½�0½�½�½P   P   ��������E���f�����������:�����������z½�#½X5½�C½�M½ZQ½�M½�C½y5½�#½�½P   P   9 ½���i�������?��� �������$�������: ½�½&½X5½	A½�G½tG½@A½�5½/&½ ½P   P   ½����V�������C�������X�������@���N����½�½�#½�0½48½�:½A8½�0½�#½
½P   P   y ½��������k���������������������_���N���: ½z½�½�%½�*½�*½�%½�½�½P   P   
������~���v�����������F��������������@������������½�½�½Q½�½?½�½P   P   ����$��������������������������������������$�������W���=���Z½�½½�½h���P   P   ����H���x�������������7�������F�������X�������:�������"���U����������'���h���P   P   ����������������k�������������������������� �������R���l���w������h���Z���c���P   P   ����������w�������k�����������������C���?����������$�����������������������P   P   ����1�����������w��������������v���k�����������f���!�������|�����������V���i���P   P   �����������������������x�������~�������V���i���E����������w���������������2���P   P   b���h�������1����������H���$���������������������	���N�����������w���N���F���P   P   �����������R������;���0����������½�½�½%���������������������Գ��q���P   P   q���U�������μ�������������� ½�½�½�½�½�½�½����+���#�����������p���P   P   Գ����������������� �������	½�½%+½�4½8½�4½�*½�½`	½~���������������P   P   ���)���/��������������/����½u$½�7½�E½N½N½�E½�7½Z$½o½������������P   P   ����������������=������u½w&½?½sQ½']½~a½]½5Q½�>½j&½o½~���#���P   P   ���Q�������˿���������W���Y	½[$½?½�U½�d½8m½Pm½e½�U½�>½Z$½`	½+���P   P   ����J�������}��������������������½�7½5Q½e½or½Sw½Gr½e½5Q½�7½�½����P   P   ��������������������������������½�*½�E½�\½7m½$w½Sw½Pm½]½�E½�*½�½P   P   %�������$�����������9������a�������D½�4½�M½\a½7m½or½8m½~a½N½�4½�½P   P   �½��������I������������������I���j½T½�7½�M½�\½e½�d½']½N½8½�½P   P   �½:���0�������ۼ��Q������t������������½T½�4½�E½5Q½�U½sQ½�E½�4½�½P   P   �½M���2�������������ϵ������������������j½D½�*½�7½?½?½�7½%+½�½P   P   �������O������Ļ����������b���л����������I��������½�½[$½w&½u$½�½�½P   P   �������
�������&�������(���N���b�������t�������a�����������Y	½u½�½�	½ ½P   P   0��� �����������0�����������(�������ϵ��������������������W������/����������P   P   ;����������X������ܹ�����������������Q�������9���������������=������� �������P   P   �������[���q����������0���&���Ļ������ۼ����������������������������������P   P   R���p���2�������q���X���������������������I����������}���˿������������μ��P   P   ���x������2���[����������
���O���2���0�������$������������������/�����������P   P   ��������w���p����������� �����������M���:���������������J���Q������)�������U���P   P   ֐�������������a���#���m���	����½F½�½F½U½i���9�����������Z���0������P   P   ���ԓ��Y���������f�������½�½#'½�/½e/½'½�½�½�������������8���P   P   0���9���|�����������r������%½!+½�?½�L½Q½tL½K?½�*½�½����4���8������P   P   Z�������z���^������G�������S½66½Q½�c½�m½�m½�c½�P½6½-½����4������P   P   ��������������������������F½:½�Y½�r½��½��½U�½�r½�Y½�9½-½��������P   P   ����ù��ĭ�������������6����½�5½�Y½�w½�½ٙ½��½$�½�w½�Y½6½�½���P   P   9���0���������"���p�������½�*½�P½�r½�½W�½ɥ½3�½$�½�r½�P½�*½�½P   P   i�����������I��������������f����½�>½�c½F�½ޙ½��½ɥ½��½U�½�c½K?½�½P   P   U½����<���ٴ��b�������������½�&½BL½Mm½׈½ޙ½W�½ٙ½��½�m½tL½'½P   P   F½P�������m����������������������
½/½�P½Mm½F�½�½�½��½�m½Q½e/½P   P   �½����@������D���ݤ��q�����������H���½/½BL½�c½�r½�w½�r½�c½�L½�/½P   P   F½�������������������d���U�������0���H����
½�&½�>½�P½�Y½�Y½Q½�?½#'½P   P   �½����o���)�����������[���E���ɧ��������������½�½�*½�5½:½66½!+½�½P   P   	�����������)���ި������ۖ�����E���U���������������f����½�½F½S½%½½P   P   m���C�����������Ǫ������Ҙ��ۖ��[���d���q����������������6������������������P   P   #���
������S������v�������������������ݤ�������������p����������G���r���f���P   P   a����������²��,������Ǫ��ި����������D������b������"��������������������P   P   ����Ϋ��U�������²��S�������)���)���������m���ٴ��I�������������^����������P   P   ����ؠ��*���U������������������o�������@�������<����������ĭ������z���|���Y���P   P   ���]���ؠ��Ϋ�����
���C�������������������P�����������0���ù����������9���ԓ��P   P   n���r��~��,��������������������½½½�½�½����B���$��� ��������}��Vr��P   P   Vr��dr��B}��������� ���8����½�&½':½�D½OD½�9½U&½|½����������������*}��P   P   �}��x���}���������.��������½�>½�Z½[m½�r½mm½~Z½�>½N½k���������������P   P   ����S���-���Ԑ��Ϊ����������#½O½,r½��½��½��½݌½�q½�N½�#½n�����������P   P    ������ ������%�������{����#½U½�~½1�½9�½@�½�½5�½�~½�T½�#½k�������P   P   $���¤��K���Y������� �������a½�N½�~½;�½��½p�½��½��½��½�~½�N½N½����P   P   B���<���9���Ϙ��3���^������H½|>½�q½�½��½��½D�½z�½��½5�½�q½�>½|½P   P   ��������Ϋ��2���&���������������"&½>Z½̌½�½j�½�½D�½��½�½݌½~Z½U&½P   P   �½����Z�������җ������2���>���>½�9½ m½7�½9�½j�½��½p�½@�½��½mm½�9½P   P   �½X����������W���2���k���߾�������½D½wr½7�½�½��½��½9�½��½�r½OD½P   P   ½�����������x���(���j�������@���r����½D½ m½̌½�½;�½1�½��½[m½�D½P   P   ½������������������r�����������=���r����½�9½>Z½�q½�~½�~½,r½�Z½':½P   P   �½��������(���2���^~���x��~����������@�������>½"&½|>½�N½U½O½�>½�&½P   P   ������������9���9���Y~���v���v��~����������߾��>�������H½a½�#½�#½�½�½P   P   ����i�������!������Ԃ��_y���v���x��r���j���k���2��������������{�����������8���P   P   �������i���J���֓������Ԃ��Y~��^~������(���2�����������^��� ����������.��� ���P   P   ����[���Ƞ��؜������֓�����9���2������x���W���җ��&���3�������%���Ϊ���������P   P   ,���O����������؜��J���!���9���(�����������������2���Ϙ��Y������Ԑ���������P   P   ~������ϋ�����Ƞ��i��������������������������Z���Ϋ��9���K��� ���-����}��B}��P   P   �r��Ex������O���[������i�������������������X�����������<���¤�����S���x��dr��P   P   �?���E���U���n��Ύ�������������C½!!½'½� ½½����I���#���0���bn��CU��ME��P   P   ME���E���R��}m��V�������c����½:½VU½�b½rb½�T½�9½)½������������m��fR��P   P   CU���M��pU��[m��J�������u����+½[½À½�½7�½Ԙ½u�½�Z½P+½���� ������m��P   P   bn��p\��Z\���n���������3����6½p½�½t�½��½��½L�½��½�o½e6½���� �������P   P   0���1q���f��kq�����)�������6½�v½��½�½��½	ý��½��½��½rv½e6½��������P   P   #��������t��ot������R�������p+½�o½��½��½ý0(ý?(ýý��½��½�o½P+½����P   P   I���,��������x��߃��������½pZ½��½��½ýO3ý�>ý23ýý��½��½�Z½)½P   P   �������������}���}������X�������Z9½P�½�½��½(ý�>ý�>ý?(ý��½L�½u�½�9½P   P   ½������������v��;���l�������u½�T½R�½t�½�ý(ýO3ý0(ý	ý��½Ԙ½�T½P   P   � ½����2�������br��ur����������)���i ½�a½Π½t�½��½ýý��½��½7�½rb½P   P   '½�������_���n��Ee���m���������+���?&½�a½R�½�½��½��½�½t�½�½�b½P   P   !!½�������]����k��s[��][��|k�����?���+���i ½�T½P�½��½��½��½�½À½VU½P   P   C½������������k���U��]O���U��k���������)���u½Z9½pZ½�o½�v½p½[½:½P   P   �����������������k��V��hJ��0J���U��|k�����������������½p+½�6½�6½�+½�½P   P   ����N���2���N����n���[���O��hJ��]O��][���m������l���X�������������3���u���c���P   P   ���ߤ������o���>s���e���[��V���U��s[��Ee��ur��;����������R���)��������������P   P   Ύ������΄���~���w��>s���n���k���k���k��n��br���v���}��߃�������������J���V���P   P   �n���q��9u���y���~��o���N�����������]���_������������}���x��ot��kq���n��[m��}m��P   P   �U���\���g��9u��΄������2�����������������2����������������t���f��Z\��pU���R��P   P   �E��KN���\���q������ߤ��N�����������������������������,�������1q��p\���M���E��P   P   ���<	������A���l�����$��������½2½�8½�1½½X���%������?l��A��������P   P   ���0	�����&?���p��`�������1"½�S½Ex½݋½��½�w½�R½~!½���������o���>����P   P   ��������?��pq��a������-@½�½��½h�½��½�½`�½k�½�?½����Ȱ��4q���>��P   P   A��%'��/'��YA��p��C�������P½Q�½��½�ý�)ý~)ý^ýR�½֜½\P½����Ȱ���o��P   P   ?l��gC��6���C��l��ҩ�������P½��½T�½�6ý�_ý�mý�_ýG6ý�½��½\P½��������P   P   ����d���H���H���d��,��������?½�½;�½Cý�{ýQ�ý�ý�{ý8Cý�½֜½�?½����P   P   %���4���x]���M��S]���������!½�½"�½E6ý�{ýa�ý��ý��ý�{ýG6ýR�½k�½~!½P   P   X���E���@r���T���T��Fr����������R½<�½�ý�_ý�ý��ý��ý�ý�_ý^ý`�½�R½P   P   ½�������4[���L���Z��?��������½tw½~�½))ý:mý�ýa�ýQ�ý�mý~)ý�½�w½P   P   �1½��������`���E���E���`��]���B����0½*�½5�½))ý�_ý�{ý�{ý�_ý�)ý��½��½P   P   �8½&���/���e���@��3���?���d������H���18½*�½~�½�ýE6ýCý�6ý�ýh�½݋½P   P   2½Q���,����g���<��M%��B%���<���f��;���H����0½tw½<�½"�½;�½T�½��½��½Ex½P   P   �½8���y����g���;�����8��~���:���f������B����½�R½�½�½��½Q�½�½�S½P   P   �����������f��%=�����{����~���<���d��]������������!½�?½�P½�P½-@½1"½P   P   $���Y���H����a��A��&��`��{��8��B%���?���`��?���������������������������P   P   �������s��4\���F���3��&��������M%��3���E���Z��Fr�����,���ҩ��C���a���`���P   P   �l���e���^���U���M���F��A��%=���;���<���@���E���L���T��S]���d��l��p��pq���p��P   P   �A���D���I��O���U��4\���a��f���g���g��e���`��4[���T���M���H���C��YA��?��&?��P   P   ����'���6���I���^���s��H�������y���,���/����������@r��x]���H��6��/'�������P   P   <	��S���'���D���e�����Y������8���P���&����������E���3����d��gC��%'�����0	��P   P   B�������E������=��/~��Y���i���6+½tJ½&T½�I½l*½��������|��H<�����z���3���P   P   3���x������� ��`C���������-4½�w½�½��½��½��½ w½'3½����א��B�� ������P   P   z������������ ���D��T��������\½��½-�½z(ý8ý�'ý��½��½�[½�������D�� ��P   P   �����������5���B�����z½�q½��½\6ý�xý#�ý!�ý�xý�5ýh�½�p½�½���B��P   P   H<��i���������@<��;�������5q½��½vVýW�ý�ý��ý.�ý�ýVýO�½�p½���א��P   P   �|���3��M��0���3���|������\½��½PVý��ýM
Ľ�1Ľ=1Ľ
Ľ��ýVýh�½�[½����P   P   ����c���)��{��`)��]c��+���:3½Գ½�5ý
�ý
Ľ�EĽ�[ĽhFĽ
Ľ�ý�5ý��½'3½P   P   ��������RE��������XE���������rv½��½xý��ýR1Ľ�[Ľ�[Ľ=1Ľ.�ý�xý��½ w½P   P   l*½ո���_���&��l��&��_��L���*½��½U'ý��ý��ýR1Ľ�EĽ�1Ľ��ý!�ý�'ý��½P   P   �I½�����t���-��Q��l���-���s�������H½��½17ý��ý��ý
ĽM
Ľ�ý#�ý8ý��½P   P   &T½����Q���G4��v����������3����������[S½��½U'ýxý
�ý��ýW�ý�xýz(ý��½P   P   tJ½���2���~7����������l���d����6����������H½��½��½�5ýPVývVý\6ý-�½�½P   P   6+½���т���7������1��������������6����������*½rv½Գ½��½��½��½��½�w½P   P   i�������u��
5��S�������-�����������d����3���s��L������:3½\½5q½�q½�\½-4½P   P   Y�������`��/��J��r���O���-������l�������-��_������+�����������z½��������P   P   /~���d���F���'���	������r�������1�����������l��&��XE��]c���|��;������T������P   P   =��5���*��Y������	��J��S�����������v��Q��l�����`)���3��@<���B���D��`C��P   P   �����������Y���'��/��
5���7��~7��G4���-���&�����{��0�����5��� ��� ��P   P   E��������������*���F���`���u��т��2���Q����t���_��RE���)��M�����������������P   P   ����,����������5���d����������������������ո�������c���3��i����������x���P   P   �<���J���q�����B����V��!��������@½�i½�x½Mi½�?½���������T�����������p��J��P   P   J��PJ���k������F��p������K½�½��½�ý�ý�½�½sJ½�����n�����ë��k��P   P   �p��@]���p����������}��� ½
�½M�½7Zý1�ý�ýޗý�YýS�½��½a���||����ë��P   P   ����H�������������=}��T½N�½�1ý�ý�Ľ%5Ľ
5Ľ>Ľ�ý�0ý|�½�
½||�����P   P   ����д������Դ������Bo�� ½�½uBý�ý]LĽ0�Ľ�Ľ&�ĽHLĽ��ý�Aý|�½a����n��P   P   �T������U���K������U������$�½�0ý��ýeĽ��Ľ�Ž�Žn�Ľ@eĽ��ý�0ý��½����P   P   ����`2��X�������O���2������gJ½a�½�ýLĽZ�ĽeŽ�<Ž�Žn�ĽHLĽ�ýS�½sJ½P   P   ����_p��N����������2�� p�����l�½+Yý�ĽїĽ�Ž�<Ž�<Ž�Ž&�Ľ>Ľ�Yý�½P   P   �?½U����,��������������S,������?½p�½�ýp4Ľc�Ľ�ŽeŽ�Ž�Ľ
5Ľޗý�½P   P   Mi½����SI��3����������������H�������g½�ýԫýp4ĽїĽZ�Ľ��Ľ0�Ľ%5Ľ�ý�ýP   P   �x½����\����������&���J��������Z������qw½�ý�ý�ĽLĽeĽ]LĽ�Ľ1�ý�ýP   P   �i½(����b�����֧��4���~��7�������9a�������g½p�½+Yý�ý��ý�ý�ý7Zý��½P   P   �@½�����\��;���:���Ps��Ga���r����������Z������?½l�½a�½�0ýuBý�1ýM�½�½P   P   ���������J��V��������s��!X���W���r��7��������H���������gJ½$�½�½O�½
�½�K½P   P   "����q��A.�������������a��!X��Ga���~��J�������S,�� p���������� ½T½� ½���P   P   �V��4��+
������e���}�������s��Ps��4��&�����������2��2��U��Bo��=}���}��p��P   P   B�������1�����������e����������:���֧������������������O����������������F��P   P   ���N���(�������������������V���;����������3���������������K���Դ�������������P   P   �q������R���(���1���+
��A.���J���\���b��\��SI���,��N��X���U������������p���k��P   P   �J��^������N�������4���q����������(�����������U���_p��`2������д��H���@]��PJ��P   P   ��������j쿽�?��X���# ��?���n½�\½��½Ũ½E�½�[½�½.���������	>��j뿽����P   P   ����R���?俽y;�������B������.m½�½�Eý�vý1vý�Dý��½�k½����:A��:���$:��8㿽P   P   j뿽�Ͽ��뿽;��6���nU���½�½�Zý��ýi1ĽNĽ+1Ľ�ý}Yý��½�½�S��ص��$:��P   P   	>��H ��� ���>������T��U½J�½�ýeLĽ�Ľ�ŽYŽT�Ľ{KĽ!�ýA�½`½�S��:���P   P   ����rE��8$��wE�������A���½0�½7�ý˅Ľ�'Žw�Ž��Ž;�Žs'ŽJ�Ľ<�ýA�½�½:A��P   P   ������xP���P��+���Q������½�ý��ĽjHŽ��ŽZ"ƽ]"ƽ��Ž�GŽJ�Ľ!�ý��½����P   P   .�����������^����������2���kk½�Yý�KĽ"'Ž��Ž�Hƽ~nƽ�Hƽ��Žt'Ž{KĽ}Yý�k½P   P   �½B��g����n��@n��%���2B��1½/�½=�ý��Ľ�Ž"ƽdnƽ~nƽ]"ƽ;�ŽT�Ľ�ý��½P   P   �[½�������a~���Y��3~���������Z½�CýB0Ľ�Že�Ž"ƽ�HƽZ"ƽ��ŽYŽ+1Ľ�DýP   P   E�½9����������I���I��:���:�������½�tý�LĽ�Ž�Ž��Ž��Žw�Ž�ŽNĽ1výP   P   Ũ½_���.(�� ���/=��2���<������&�������½�týB0Ľ��Ľ"'ŽjHŽ�'Ž�Ľi1Ľ�výP   P   ��½�����0������6���������M5��.���/��������½�Cý=�ý�KĽ��Ľ˅ĽeLĽ��ý�EýP   P   �\½R����(�����P3���/ֿ����1��.����&������Z½/�½�Yý�ý7�ý�ý�Zý�½P   P   n½����������7����ȿ��ȿ���M5�����:�����1½kk½�½0�½J�½�½.m½P   P   @����D�����������>������T׿��ȿ�/ֿ�����<��:������2B��2�������½U½�½����P   P   # ���������Ԁ���K��%������������2���I��3~��%�������Q���A���T��nU���B��P   P   X���0�������p��\���K���>��7��P3��6��/=���I���Y��@n������+����������6�������P   P   �?��+G���R��`a���p��Ԁ���������������� ������a~���n���^���P��wE���>��;��y;��P   P   j쿽��a&���R�����������������(���0��.(���������g������xP��8$��� ���뿽?俽P   P   �����п���+G��0�������D������R�������_���9������B����������rE��H ���Ͽ�R���P   P   ؾ�z��7��o���6�������w��H½��½5�½�½��½�½�	½%u��a���3�����^6���ﾽP   P   �ﾽ	�-��!����D�����g�����½�Cýg�ý�ĽKĽ�ý9Býɗ½����g���B��O����+��P   P   ^6������6��d����I������½� ý��ý+�ĽQŽs)Ž�Ž�Ľ��ý��½n½o���G��O���P   P   ����S���S��ץ���C�����K"½7ýaAĽ�&Ž��Ž)ƽ�(ƽ��Ž�%Ž�?Ľ�5ý� ½o���B��P   P   3������ہ��访��3��1��m½�6ý�dĽ�wŽyTƽ��ƽ�ǽ0�ƽ�SƽwŽ�cĽ�5ýn½g��P   P   a���u������/����������}���U�½%@Ľ�wŽ��ƽ�Eǽ�ǽ#�ǽ�Eǽ��ƽwŽ�?Ľ��½����P   P   %u������|��]ο����}���u����½+�ý&Ž�SƽqEǽ��ǽ�ȽV�ǽ�Eǽ�Sƽ�%Ž��ýɗ½P   P   �	½.��?H���俽b俽�G�����	½�Aý�Ľ(�Ž��ƽ��ǽ�Ƚ�Ƚ#�ǽ0�ƽ��Ž�Ľ9BýP   P   �½�g��Ȉ��\���?ʿ�7�������zf��݀½��ý� Ž�'ƽǽ��ǽ��ǽ�ǽ�ǽ�(ƽ�Ž�ýP   P   ��½��������������\������ʼ��������½� Ľ�'Ž�'ƽ��ƽqEǽ�Eǽ��ƽ)ƽs)ŽKĽP   P   �½:�������# ��?����y�������������W�����½� Ľ� Ž(�Ž�Sƽ��ƽyTƽ��ŽQŽ�ĽP   P   5�½��������(�� ����P��^P���'������W�����½��ý�Ľ&Ž�wŽ�wŽ�&Ž+�Ľg�ýP   P   ��½����\���7)��㗿�a;�����m:�����'����������݀½�Aý+�ý%@Ľ�dĽaAĽ��ý�CýP   P   H½�i�������!��6����;��l	��	��m:������ʼ��zf��	½��½U�½�6ý7ý� ý��½P   P   �w�����`���*�����0R�����l	�����^P����������������u��}���m½K"½�½g���P   P   ����u���.K��_���H���5|��0R���;��a;���P���y��\���7����G��}�������1�����������P   P   6��Q ������翽|Ϳ�G������6���㗿� ���?�������?ʿ�b俽�������3���C���I���D��P   P   o���������gѿ��翽_���*���!��7)���(��# �����\����俽]ο�/���访�ץ��d���!���P   P   �7���U������������.K��`�������\���������������Ȉ��?H��|������ہ���S���6��-��P   P   z�m���U�����Q ��t�������i���������:�������g��.������u�������S�����	�P   P   �Ľ��彽�D��۾������q��(N��½��½)#ýxFý2"ýn�½%½�J��	n��	���ؾ��B���佽P   P   �佽%彽�7���Ծ�Ů������������½��ý�jĽr�Ľ��Ľ!iĽR�ý��½�����������vҾ�6��P   P   �B�����C���Ӿ�2�������s½rdý��ĽF�Ž�#ƽ�Zƽ�"ƽ��Ž��Ľ�aý�½1������vҾ�P   P   ؾ��i��j��پ�����/���5½��ý@Ž�Uƽx=ǽ�ǽ��ǽ�<ǽvTƽPŽ��ý�2½1������P   P   	����㾽���/侽��������"½0�ý�IŽD�ƽ��ǽ��Ƚ?�Ƚ-�Ƚ��ǽ�ƽHŽ��ý�½����P   P   	n��gw��-���v����w���n�������bý�Ž��ƽ4ȽyBɽ��ɽg�ɽ8Bɽ�3Ƚ�ƽPŽ�aý����P   P   �J��U���Q��V���Q��x���J����½��Ľ�Tƽ��ǽ1BɽMʽ!fʽGʽ8Bɽ��ǽvTƽ��Ľ��½P   P   %½����ׯ���+��{+������$����½��ý��Ž�;ǽ¹Ƚ�ɽ�eʽ!fʽg�ɽ-�Ƚ�<ǽ��ŽR�ýP   P   n�½�6���	���I�����cI�����q5���½�gĽ�!ƽo�ǽ'�Ƚ�ɽMʽ��ɽ@�Ƚ��ǽ�"ƽ!iĽP   P   2"ýߙ���R��g���뾽5뾽f���Q������) ý��Ľ�Xƽo�ǽ¹Ƚ1BɽyBɽ��Ƚ�ǽ�Zƽ��ĽP   P   xFý�������}���־������վ�u{�����o����Cý��Ľ�!ƽ�;ǽ��ǽ4Ƚ��ǽx=ǽ�#ƽr�ĽP   P   )#ý����z������6ʾ��f��bf���Ⱦ�ɇ������o���) ý�gĽ��Ž�Tƽ��ƽD�ƽ�UƽF�Ž�jĽP   P   ��½������������Ǿ�.K�����J���ž�ɇ����������½��ý��Ľ�Ž�IŽ@Ž��Ľ��ýP   P   ½+9��8U��
���˾��K�����&��J���Ⱦ�u{���Q��q5���½��½�bý0�ý��ýrdý��½P   P   (N�����B��j���ؾ��h��� ��������bf���վ�f�����$����J������"½5½s½����P   P   �q��$������MM��������h���K��.K���f������5뾽cI������x���n������/�����������P   P   ����5{���U���/�������ؾ��˾��Ǿ�6ʾ��־��뾽���{+���Q���w����������2���Ʈ��P   P   ۾�羽���R���/��MM��j��
���������}��g���I���+��V��v���/侽پ��Ӿ��Ծ�P   P   �D��kl����������U������B��8U�����z�������R���	��ׯ���Q��-������j���C���7��P   P   �彽��kl��羽5{��$�����+9��������������ߙ���6������U��gw���㾽�i����%彽P   P   ,T������<���iǽ��Ǿ�}뿽@��p'½�ý��ýu�ý�ý�ý�#½����濽�þ��ý��������P   P   ������������%徽[E�����/-ý�kĽ�UŽJ�Ž��Ž�SŽ�hĽ:)ý���A��K᾽����켽P   P   ����Ի����������$ﾽu���,½��ý��Ž��ƽO�ǽY Ƚ�ǽ��ƽŽ!�ý@)½�q��e쾽����P   P   �ý�_/���/���Ľ��㾽Pt���R½UĽ�Iƽo�ǽC;ɽ3�ɽ��ɽ�9ɽC�ǽ#GƽRĽ�O½�q��K᾽P   P   �þ��ҽ�d���oӽ��ľ��B��9+½+TĽ�ƽ)�Ƚ�7ʽ�I˽��˽;I˽�6ʽK�Ƚ�ƽRĽ@)½A��P   P   �濽Ȗ���齽�齽L����翽3���R�ýuHƽ]�ȽϏʽD̽��̽m�̽�̽�ʽK�Ƚ#Gƽ!�ý���P   P   ����m���c��"	���c���m�����q)ý։ŽY�ǽ�6ʽ�̽�5ͽa�ͽ6ͽ�̽�6ʽC�ǽŽ:)ýP   P   �#½�>��L徽�/���/�� 徽`>��#½+hĽ��ƽ 9ɽ�H˽�̽_�ͽa�ͽm�̽;I˽�9ɽ��ƽ�hĽP   P   �ýg����]��;Z��^���Y���\��A���1ý�QŽ=�ǽF�ɽ˧˽�̽�5ͽ��̽��˽��ɽ�ǽ�SŽP   P   �ý�~��(���ʁ���۽�F۽�����.���m|����ý��Ž��ǽF�ɽ�H˽�̽D̽�I˽3�ɽY Ƚ��ŽP   P   u�ý����6��ڡ���½�u������
���� ��I�����ý��Ž=�ǽ 9ɽ�6ʽϏʽ�7ʽC;ɽO�ǽJ�ŽP   P   ��ý5���(��o���󳽽�-��-������|������I�����ý�QŽ��ƽY�ǽ]�Ƚ*�Ƚo�ǽ��ƽ�UŽP   P   �ý�����1����������lϼ����S���|���� ��m|��1ý+hĽ։ŽuHƽ�ƽ�Iƽ��Ž�kĽP   P   q'½����Ŀ�E���m���
��
��� ����������
���.���A���#½q)ýR�ý+TĽUĽ��ý/-ýP   P   @��uC���a�������Ž�0���м�
���lϼ�-�����������\��`>�����3���9+½�R½�,½���P   P   }뿽qr��?꾽�^��ཽ�x��0��
������-��u��F۽��Y�� 徽�m���翽�B��Pt��u��[E��P   P   �Ǿ�����i��5��w��ཽ�Ž�m�������󳽽�½��۽�^���/���c��L����ľ��㾽%ﾽ&徽P   P   iǽ�>׽��_��5���^������E���0���o���١��ʁ��;Z���/��"	���齽oӽ��Ľ���������P   P   <����2��v����i��?꾽�a��Ŀ���(��6��(����]��L徽�c���齽d����/��������P   P   ���� ����2��>׽�����qr��uC���������5��������~��g����>���m��Ȗ���ҽ�_/��Ի�����P   P   5i��[���pL���W��-����7��!����@½1qý�6Ľ�{Ľw4Ľ�mý,<½F���z1��ɩ���R���H������P   P   ����J����4���N���ؽ�ֲ��������ýR\Ž�ƽJǽ#Iǽ��ƽXŽ<�ýʭ��-���ӽ��J��=2��P   P   �H��[�nJ���M��S潽c����I½q�Ľ��ƽ�Ƚ�ɽ/Kʽ��ɽ�Ƚ(�ƽ��Ľ�D½��x⽽�J��P   P   �R�����������T��Zֽ���N½d>ŽP�ǽ�Dʽ�̽l�̽��̽��˽�Aʽ��ǽF:Ž?{½��ӽ�P   P   ɩ���c������d��{��������G½=ŽiGȽ�˽ybͽ�νLfϽ)�ν�`ͽ˽�DȽF:Ž�D½-���P   P   z1���l��l�������]m���2��A���e�Ľ��ǽ�˽@�ͽ��Ͻ'ѽ�ѽ��Ͻ �ͽ˽��ǽ��Ľʭ��P   P   F���ꌾ�2%��W���p%��O��������ý?�ƽ"Bʽ[aͽ��Ͻ�ѽm&ҽ �ѽ��Ͻ�`ͽ�Aʽ)�ƽ<�ýP   P   ,<½�����ҽ��ݼ��ݼ�Tҽ�৿�U;½vWŽ_�Ƚ��˽9�ν\ѽ|&ҽm&ҽ�ѽ)�ν��˽�ȽXŽP   P   �mý�����w�����ܠ������v�������ký#�ƽ4�ɽ��̽/eϽ\ѽ�ѽ'ѽLfϽ��̽��ɽ��ƽP   P   w4Ľ|\�� ���P��Tq���p���O��}����Y���1Ľ�Eǽ<Hʽ��̽9�ν��Ͻ��Ͻ�νl�̽/Kʽ#IǽP   P   �{ĽH����Z���}���P���绽iO���{���W�����KwĽ�Eǽ4�ɽ��˽[aͽ@�ͽzbͽ�̽�ɽJǽP   P   �6Ľ����{��$����>������I���1<�������v������1Ľ#�ƽ_�Ƚ"Bʽ�˽�˽�Dʽ�Ƚ�ƽP   P   1qýj_��]��6����8��VZ��=���X���5�������W���Y���kývWŽ?�ƽ��ǽiGȽP�ǽ��ƽR\ŽP   P   �@½֧���������U@���[��&庽亽�X��1<���{��}�������U;½�ýe�Ľ=Žd>Žr�Ľ��ýP   P   !���<���}���U���T��������&庽=��I���iO���O���v��৿�����A����G½N½�I½����P   P   �7��/���
ٽ�����v���뻽����[��VZ�������绽�p�����Tҽ�O����2��������c���ֲ��P   P   -����r���+��C伽"����v���T��U@���8���>���P��Tq��ܠ���ݼ�p%��]m��{���Zֽ�S潽�ؽ�P   P   �W���i����������C伽����U������6���$����}���P������ݼ�W��������d���T���M���N��P   P   pL���������������+��
ٽ�}�����]��{���Z�� ���w���ҽ�2%��l����������nJ���4��P   P   [�����������i���r��/���<���֧��j_������H���|\����������ꌾ��l���c������[�J���P   P   Iݷ��)��~
��>m��l9��SI���l��/j½g	ĽaŽFxŽ�Ž�Ľ�c½�d��WA��B2��(g�����L'��P   P   L'��W(���븽�c��t����������TĽ��ƽYiȽBVɽUɽ�eȽ�ƽNĽ�����쾽�m���^���踽P   P   �����������b�������M���z½��ŽY�Ƚ�O˽�̽,�ͽ�̽�K˽6�Ƚ=�Ž�s½�G������^��P   P   (g���[���\��i���q���L����½Y�ƽ�8ʽzͽR�Ͻ�0ѽ�/ѽ��Ͻvͽb3ʽ�ƽ��½�G���m��P   P   B2���{��D繽�|���4���x½��ƽl�ʽ?�ν��ѽ��ӽi�ԽQ�ӽ��ѽ��ν��ʽ�ƽ�s½�쾽P   P   WA��aܻ�ӟ��'���lݻ�*C������ؾŽ�6ʽ՟νӀҽ:gս��ֽ��ֽ�eս,ҽ��νb3ʽ=�Ž����P   P   �d��`��{z���ֺ��z���`���e��?OĽ��Ƚ�vͽ�ѽ�fս+�׽ �ؽ¿׽�eս��ѽvͽ6�ȽNĽP   P   �c½�᾽�c��������&c��*᾽�b½r�ƽ#K˽�ϽR�ӽ�ֽߑؽ �ؽ��ֽQ�ӽ��Ͻ�K˽�ƽP   P   �Ľ�5��fD��fk���ɺ��j��BC��$4��{Ľ7cȽP�̽:-ѽ"�Խ�ֽ+�׽��ֽi�Խ�/ѽ�̽�eȽP   P   �Žy4��& ��u���f���݋��и��'���1���Ž�Pɽzͽ:-ѽR�ӽ�fս:gս��ӽ�0ѽ,�ͽUɽP   P   FxŽ����}��g����d���ڹ��b������y��r����rŽ�PɽP�̽�Ͻ�ѽӀҽ��ѽR�Ͻ�̽BVɽP   P   aŽ����:�������N��7_��V^���K��f������r����Ž8cȽ#K˽�vͽ՟ν@�νzͽ�O˽YiȽP   P   g	Ľ`8�����'���I��� ��G�������E��f��y��1��{Ľr�ƽ��Ƚ�6ʽl�ʽ�8ʽY�Ƚ��ƽP   P   /j½�;�����C����P��L"������u�������K������'���$4���b½?OĽؾŽ��ƽZ�ƽ��Ž�TĽP   P   �l�� 龽 K��^���i���b��{�������G���V^���b��и��BC��*᾽�e������x½��½�z½����P   P   SI��&h���k���r�����F๽�b��L"��� ��7_���ڹ�݋���j��&c���`��*C��𾽔L���M�����P   P   m9��F份܂���$���Ѻ����i���P���I���N���d��f����ɺ�����z��lݻ��4���q������t��P   P   >m��"�������ߺ��$���r��^���C���'�����g���u���fk������ֺ�'����|��i���b���c��P   P   ~
���a��������܂���k�� K��������:���}��& ��fD���c��{z��ӟ��D繽�\������븽P   P   �)������a��"���F份&h�� 龽�;��`8����������y4���5���᾽`��aܻ��{���[������W(��P   P   �����贽���緽�L�����a�w�½%�Ľ�Yƽi�ƽpVƽ��Ľ֟½�追���C��(߷��
���崽P   P   �崽(紽�鵽X۷�q�����������GŽ�ȽR�ʽ�/̽o.̽��ʽ�xȽ�>ŽA���e�����Է��嵽P   P   �
��po�����ڷ�͹���t���½@ǽ�x˽��ν8ѽ2ҽ�4ѽ��νq˽e7ǽ^�½�l�������Է�P   P   (߷��z���{��^ⷽ왺�Ns���%ý�MȽmͽg�ѽz]սE1׽�/׽Zս��ѽ�eͽ�EȽ�ý�l������P   P   C�������0�������F��7���½�KȽ�ν��ӽiؽ۽� ܽ�۽cؽ��ӽ�ν�EȽ^�½eP   P   ���2͹�F$���$���ι�@������A;ǽ&jͽ �ӽcٽ�.ݽ�f߽Ef߽�,ݽ�ٽ��ӽ�eͽe7ǽA���P   P   �追Ի�PG��i���G��Gջ�꿽�@Ž�r˽-�ѽؽ�-ݽ���B�����,ݽcؽ��ѽq˽�>ŽP   P   ֟½�ڽ�p���nǸ�RǸ�5����ڽ�R�½�wȽ#�ν8Yս۽�e߽��B��Ef߽�۽Zս��ν�xȽP   P   ��Ľ��������+6���\���5��8�������R�Ľ��ʽ 2ѽ�,׽ܽ�e߽��འf߽� ܽ�/׽�4ѽ��ʽP   P   pVƽ\��P���򡹽����������,���7���Qƽ)̽v�ѽ�,׽۽�-ݽ�.ݽ۽E1׽2ҽo.̽P   P   i�ƽ���vZ�������ܷ�L%��۷�S���lU��ݼ����ƽ)̽ 2ѽ8Yսؽcٽjؽz]ս8ѽ�/̽P   P   �Yƽ�������Q,��P÷�������뿷�'��d���ݼ���Qƽ��ʽ#�ν-�ѽ �ӽ��ӽg�ѽ��νR�ʽP   P   %�ĽX���]��.������3��?���1��U���'��lU��7��R�Ľ�wȽ�r˽&jͽ�νmͽ�x˽�ȽP   P   w�½!���z�������hƷ�I5��-f���d��1��뿷�S���,�������R�½�@ŽA;ǽ�KȽ�MȽ@ǽ�GŽP   P   a�,佽^���c����ⷽ����+���-f��?������۷�����8����ڽ�꿽������½�%ý�½����P   P   ����޻�l���y?������,������I5���3�����L%������5��5���Gջ�@��7�Ns���t�����P   P   �L��V׹��Q���Ѹ��f������ⷽhƷ����P÷��ܷ�����\��RǸ��G���ι��F��왺�͹��q���P   P   緽5��@.��fs���Ѹ�y?��c�������.��Q,������򡹽+6��nǸ�i���$������^ⷽڷ�X۷�P   P   �������9��@.���Q��l���^���z����]�����vZ��P�������p���PG��F$���0���{������鵽P   P   �贽�s������4��V׹��޻�,佽!���X���������\�������ڽ�Ի�2͹������z��po��(紽P   P   '�������.������ŷ�4t��sU��OýYƽRȽ��Ƚ'Ƚ�ƽ��½�H��Ag����������	'��̧��P   P   ̧����������O���)3��1������E�ƽi˽�]ν*н�'нXWνA�ʽ�ƽ�������>(��׃��c���P   P   	'���Z���*��d���@Z���Z���.ýSɽb(Ͻ��ӽ5׽dSؽ�0׽��ӽ�ϽXGɽ�"ý�O���P��׃��P   P   �������d���򓴽/��^X��^�ý��ʽ��ѽ�Aؽ/ݽ��߽7�߽,ݽ�9ؽ��ѽ�ʽѬý�O��>(��P   P   �������¢��}���I���X����*ý��ʽ��ҽ#�ڽ��ཨG���潄D� ����ڽ��ҽ�ʽ�"ý����P   P   Ag�����xⴽ�㴽'��k��2���Mɽs�ѽL�ڽ/^�?N轷����뽥K轻Y���ڽ��ѽXGɽ���P   P   �H��ɹ�c���<���c��˹�K��'�ƽ� Ͻq<ؽU��'M��0��/�K� ���9ؽ�Ͻ�ƽP   P   ��½o���������������������½��ʽa�ӽ�ݽ�C�\�������뽄D�,ݽ��ӽA�ʽP   P   �ƽ���������K��.��K������:�
ƽ�SνI-׽��߽G��\���0������7�߽�0׽XWνP   P   'ȽX��������ල�˴��ʴ�p޶�v�>���C
Ƚh!нIMؽ��߽�C�'M�?N轨G���߽dSؽ�'нP   P   ��Ƚk���Eݻ�S[���������ߋ��W��E׻�����Y�Ƚh!нI-׽�ݽU��/^⽥��/ݽ5׽*нP   P   RȽ����.2��&����o��4̲��ʲ��k�������)������C
Ƚ�Sνa�ӽq<ؽM�ڽ#�ڽ�Aؽ��ӽ�]νP   P   Yƽ����qỽ���vf���d��Ѵ��ia���`������E׻�>���
ƽ��ʽ� Ͻs�ѽ��ҽ��ѽb(Ͻi˽P   P   Oý��������Da��t��yf���X��(W��ia���k��W��v�:���½'�ƽMɽ��ʽ��ʽSɽE�ƽP   P   sU��o�������궽����Ѳ�~����X��Ѵ���ʲ�ߋ��p޶���������K��2����*ý^�ý�.ý���P   P   4t���ֹ�c��W���մ�����Ѳ�yf���d��4̲�����ʴ�K�����˹�k��Y���^X���Z��2���P   P   ŷ��#��p���ĵ�j:���մ����t��vf���o�������˴�.������c��'��I���/��@Z��)3��P   P   ����������I���ĵ�W��궽Da�����&���S[���ල�K������<���㴽}���򓴽d���O���P   P   �.����������p��c����������qỽ.2��Eݻ������������c��xⴽ¢��d����*������P   P   �����`����������#���ֹ�o���������������k���X�������o���ɹ�����������Z������P   P   K��� 5��K'���K��,u���W�����9�ý��ǽ�rʽ�i˽mʽ{�ǽAuývy���F���d���>�����=0��P   P   =0���2��e謽Z?�����x�������lȽ��ν�'ӽ�ս�ս2ӽ wν3]ȽD���򺽼���"4��[ᬽP   P   ���M��o"���<���?���黽��ý�*̽CԽS۽Й߽\0�,�߽�۽�4Խ�̽��ý�ڻ��3��"4��P   P   �>���խ��׭��D����绽{�Ľ�1νyؽl�M����&�뽶���Ὦؽ#νOrĽ�ڻ�����P   P   �d��a^������a��mk��3�����ýL/ν�rٽd�ܨ�N��������Ӡ�Y佃fٽ#ν��ý�P   P   �F��������b���~����L�����_#̽�ؽ�a�{�ｱX�����F���T����｡Y佮ؽ�̽D���P   P   vy��E��"���������>��}��haȽ�9Խ��[��W������������T��Ӡ��὆4Խ3]ȽP   P   Auý����
´�縱����S´�C���CvýGwν�۽��罌�����J���F������罙۽ wνP   P   {�ǽ���wⶽ�~�����*~��ᶽw��u�ǽgӽ͏߽��t���������������&��-�߽2ӽP   P   mʽR���`���9K������剰��H��p���i����eʽ/�սo(��뽌��W���X��N�����]0��սP   P   �i˽����|빽��+C��y�� A���볽q乽���� _˽/�սΏ߽���[��{��ܨ�M�љ߽�սP   P   �rʽ�����\���O��� ������(��� ���G��lR�������eʽgӽ�۽���a�d�m�T۽�'ӽP   P   ��ǽX������Q������|��ʙ��y������G��q乽i���u�ǽGwν�9Խ�ؽ�rٽzؽCԽ��νP   P   9�ý�����������%��	���"��+!��y�� ���볽p���w��CvýhaȽ_#̽L/ν�1ν�*̽�lȽP   P   ����κ�F�V��pL��A��a����"��ʙ��(��� A���H��ᶽC���}�������ý{�Ľ��ý����P   P   �W��d-���Ѵ��D�����A��	���|������y��剰�*~��S´�?���L��3���绽�黽x��P   P   ,u������i����ȱ����D���pL���%������ ��+C����������������~���nk�����?�����P   P   �K���l�������#���ȱ��V�������Q���O����9K���~��縱���b����a���D���<��Z?��P   P   K'��᭽������i����Ѵ�F𶽎����𹽣\��|빽`���wⶽ
´�"����������׭�o"��e謽P   P    5�����᭽�l������d-���κ���W�����������Q����������E�����a^���խ�M���2��P   P   8b��|:����������!��D���3u��:+Ľ��ɽ�ͽ��ν(�ͽF�ɽ�ĽV_��Yu��"��:�������]4��P   P   ]4��k7���g��岪�ﰽ�ȸ�����!�ʽ�?ӽ�ٽ48ݽ4ݽ�ٽ.ӽ��ʽ��������ܰ�[���z^��P   P   ����3U��@�������?6������Ľ�нdE۽U�佖Y����Q�j�佈1۽��Ͻ�wĽ�J&��[���P   P   :�������b������,鰽�����Ž��ҽ��)������� ��;{���w����ҽ�yŽ��ܰ�P   P   "���̪��
��Ѫ��������	�Ľ��ҽG��K����Í�*3��������n;�܋��ҽ�wĽ���P   P   Yu���讽m�����}��{���J�Ͻ���G�f����d}�|�����`�n;�����Ͻ����P   P   V_������k���֪��è��՘��2e����ʽ9۽�~�������^a�%W�3`���������w�1۽��ʽP   P   �Ľ�d���{��9��������|��Af��Ľ�/ӽ����{�����|�W�%W�|����;{��j��.ӽP   P   F�ɽ�ɼ�L�����D�������K���Ǽ��ɽݣٽiL������0�|�^a�d}�*3�!���Q��ٽP   P   (�ͽ-��.�������
���	��;��������&��͒ͽs*ݽ����������������Í������4ݽP   P   ��νV½\��⁯���� ��k���|���S��i�����νs*ݽiL��{������f���������Y�48ݽP   P   �ͽ�	½1����e����٧��ק�3���D����䷽i���͒ͽݣٽ����~��G�K�*��V���ٽP   P   ��ɽ�7���b��0������":������5��)���D����S���&���ɽ�/ӽ9۽��H����dE۽�?ӽP   P   :+Ľ�ټ��µ�����>����<��,�������5��3���|�������Ǽ�Ľ��ʽJ�Ͻ��ҽ��ҽ�н"�ʽP   P   3u��Tx��]������PŪ�~᧽;��,�������ק�k���;���K��Af��2e��{���	�Ľ�Ž��Ľ����P   P   D���۩��n����������G,��~᧽�<��":���٧� ���	�������|��՘���}�������������ȸ�P   P   �!����������_���氫����PŪ�>�������e�������
��D�������è�����-鰽?6��ﰽP   P   �����ު�^.�����_���������������0�����ၯ�������9���֪����Ѫ��������岪�P   P   ���隧����^.������n���]���µ��b��1�\��-���L���{��k���m���
��b���@����g��P   P   |:��l^��隧��ު�����۩��Sx���ټ��7���	½V½-���ɼ��d�������讽�̪�����3U��k7��P   P   �Z���f�����ߖ��Y{��+Ѳ�Y�&�ĽJ�̽1�ѽ��ӽ��ѽr�̽�Ľ�Ի������a��􁣽Gq��._��P   P   ._��c��<!��󐣽�����˵����:ν]�ٽ���罨�罋��vvٽ<�ͽ����?���ww���~�����P   P   Gq���Ü��x��/���N�In���|Ž�#ս���n�V���u ��n����Y�m��ս�^Ž�S��uܫ��~��P   P   􁣽Z���݊��@���m���`j����ƽ�ٽ���L �������
���
�g������7f�H�ؽ?�ƽ�S��ww��P   P   �a�������^�������m��s����tŽ.ٽ�A����c�J�k��d�/
���T(�H�ؽ�^Ž?���P   P   �����ۨ��������'㨽b���J���=ս�y콧��`O��C������>�\G���7f�ս����P   P   �Ի��鮽�8��ح���;���﮽�ݻ��ͽ������/��A���!��$���!�>�/
�����m��<�ͽP   P   �ĽG;��?㪽�¥��å��媽�>����Ľ�zٽ�\�U����%��)�$��$����d�g���Y�vvٽP   P   r�̽���ꔮ�T#��誤��"��Z���*����̽+}⽘���w�
���%����!���k����
�n������P   P   ��ѽ�����Ʊ�s���$�����������%±�ː��Y�ѽ}v罿��w�
����A��C�J���
�u �����P   P   ��ӽ�½���aƩ�M���+������#���8��½ʘӽ}v罘���V��0�`O�c����W�����P   P   1�ѽ�½�����v��`��������������l��Ĳ���½Y�ѽ,}⽶\����������L ���n���P   P   K�̽F���C����z��눣�VV���흽�Q���~���l��8�ː����̽�zٽ����y콒A������]�ٽP   P   &�Ľf'���ֱ�!ѩ����0Y��h8���5���Q������#���%±�*����Ľ�ͽ=ս.ٽ�ٽ�#ս:νP   P   Z�{T������-���5��������h8���흽����������Z����>���ݻ�K����tŽ��ƽ�|Ž���P   P   +Ѳ�P��U���x8����I������0Y��VV�����+��������"���媽�﮽b���s���`j��Jn���˵�P   P   Y{������cQ���٥�������5������눣�`���M���$���誤��å��;��'㨽�m��m���N񫽜���P   P   ����-�������Ĥ��٥�x8��-���!ѩ��z���v��aƩ�s���T#���¥�ح���������@���/���󐣽P   P   ��������q�����cQ��U��������ֱ�C�����������Ʊ�ꔮ�?㪽�8�������^��݊���x��<!��P   P   �f���Μ�����-�������P��{T��f'��F����½�½�������G;���鮽�ۨ�����Z����Ü�c��P   P   ��sV���"���o������ȭ�L���"�Ž нi׽v�ٽ׽��ϽA~Ž����1��������U�����:M��P   P   :M��"R������t��j���񱱽n=����ѽ,��bl� t��5l��{U���3�ѽ���8���Uj���]�����P   P   ����������p��
�� ۳�nƽ��۽��T���j	�����a	����p�>�۽�Eƽ&������]��P   P   �U��S\���`��Lc��ɀ��nֳ�WEȽ[὿���N�������A�����St���ཇ Ƚ&���Uj��P   P   ����^j��Ϛ��kr��~��̤��Cdƽ���H �s�X] �-`+��d/�IX+��N �`��&6 ����Eƽ8���P   P   1��������͚�њ��������G+����۽����&��d�#���3���<��<���3���#�`��St��>�۽���P   P   ���� ����垽����ꞽ�è�ܙ����ѽ���<��YW ��3�I�A�[�F�6�A���3��N ����p�3�ѽP   P   A~ŽB鰽�������_������4ﰽ�Ž5����-��tY+���<���F�[�F��<�JX+�������P   P   ��Ͻܒ���[���ߞ����ߞ�\��ƒ���ϽMQ�M^	��	�`/���<�I�A���<��d/�B��a	�{U�P   P   ׽E���ŉ���Ǡ����K���Š�?���⎾��׽�\������	�tY+��3���3�-`+������6l��P   P   v�ٽM����j���c������H*�����o]���_��5����ٽ�\��M^	�-��YW �d�#�Y] �����j	�t��P   P   j׽m���=y���Q��\����[���Y��󡚽�F���h��6����׽NQ���<��'��s�N��U��cl�P   P    н�����t��|V��Q������� ȓ�w{�������F���_��⎾��Ͻ5�ὸ�񽽑���H �������,��P   P   "�Žn�������p��������!𒽾쒽w{��󡚽o]��?���ƒ���Ž��ѽ��۽��[Ὢ�۽��ѽP   P   L���#	���t���۠�5Ě�{f��Γ�!� ȓ��Y������Š�\��4ﰽݙ��H+��CdƽWEȽnƽn=��P   P   �ȭ��ۨ�ò��c���[��L:��{f����������[��H*��K���ߞ������è�����ͤ��nֳ�!۳�񱱽P   P   ���`��I��-��^ڛ�[��5Ě����Q���\������������_��ꞽ�����ʀ����j���P   P   �o��ȅ��隽�Ǜ�-��c����۠��p��|V���Q���c���Ǡ��ߞ��������њ�kr��Lc���p���t��P   P   �"��q������隽I��ò���t������t��<y���j��ŉ���[�������垽�͚�Ϛ���`�������P   P   sV���	��q��ȅ��`���ۨ�#	��n�������m���L���E���ے��A鰽 �������^j��S\������"R��P   P   ���Ơ���,��b͎�����馽�>����Ž,�ӽ�ݽ��6�ݽ��ӽS�Ž���R���BX�����r��ϕ��P   P   ϕ��曂�ު���ގ��T�������*���ֽ�R����v���~����#�\Jֽg����ū��-��������P   P   r��_����"��dڎ�`����Ů��ǽ����J�$o����(J����]X��.�ݤ�u�ƽҗ���ۛ���P   P   ���M���\�������
K�����͋ɽjg�Y9	��(��.���7���7�"�-�.�&	�_-뽇Yɽҗ���-��P   P   CX������[B��#���m���嫽�ǽ`뽿�%�l
=�Z�N�qU��N�a�<�'�$�}��_-�u�ƽ�ū�P   P   R���5і��#��.(��'ߖ��Ҧ����"��1	�-%�y�B��r\���k���k�Rc\�b�B�(�$�&	�ݤ�g���P   P   ���=~��0��>4���6��ڊ���"���bֽ�<���9=�\n\�qGt��G}�At�Rc\�a�<�.��.�\JֽP   P   S�Žd�����������H�������Ž�/��]�R�-���N�
�k�cH}��G}���k��N�#�-�^X��#�P   P   ��ӽiߴ�j&��lN��Lx��~O���(��kᴽP�ӽ����]��g�7�5jU�
�k�rGt���k�qU���7�������P   P   7�ݽ�ʼ������Ж�ಏ�Ȳ��<ϖ�Ԅ��gü��ݽ��f=�g�7���N�\n\��r\�Z�N���7�(J���P   P   ��46��ZF����~���h��P{���阽S;��%��D���]��R�-�9=�z�B�l
=��.����w�P   P   �ݽ=>�����;-�������\���Z������:!������%���ݽ�����]���.%�%��(�$o����P   P   ,�ӽ�༽�R��=2������fg���]��$b������:!��S;��gü�P�ӽ�/콑<�1	���Z9	��J��R�P   P   ��Ž� ���������I���nk���d��&a��$b�������阽Ԅ��kᴽ��Ž�bֽ"��`�kg뽤�㽖ֽP   P   �>������D���疽����h��-d���d���]���Z��P{��<ϖ��(������"������ǽ΋ɽ�ǽ�*��P   P   �馽]����6���j��ʏ��z��h��nk��fg���\���h��Ȳ��~O��H��ڊ���Ҧ��嫽����Ů�����P   P   ���h����R�����"���ʏ�����I������������~��ಏ�Lx�������6��'ߖ�m��
K��a����T��P   P   b͎�֎��C���R������j���疽���=2��;-����Ж�lN������>4��.(��#�������dڎ��ގ�P   P   �,��뱈��\���C���R���6���D�������R�����ZF������j&�����0���#��[B��\����"��ߪ��P   P   Ơ������뱈�֎�g���\������� ���༽<>��36���ʼ�iߴ�d=~��5і�����N���_���盂�P   P   6<`��c�MPn�S'��~ ��1�������Ž2 ؽ�N�`��5彾�׽XMŽ�˰�7[���Ќ�1��rn���c�P   P   ��c���c�Q-m�H��	P������佽A۽�`��{+	��Z� R�n	�� ���7۽�������9 ���%���m�P   P   rn��6h�2:n��B���&������~�ƽ^��Z�� �0�Ϯ5���/��� ��1�cc��ƽW��"����%��P   P   1����q��q�'��E�������Dʽ�������|5�R�O��]_��Q_�ӏO�qR5�Q������ ʽW��: ��P   P   �Ќ�����w����	쌽�㣽v�ƽ
�������A���g��Ƃ�)q��&���>�g��A��������ƽ����P   P   7[������Cq���v���É�5y���ɽ���&��j�A�	q�p����<���7���z��?�p��A�Q��cc����P   P   �˰�m���7���s���y���6����氽[۽�F��i5���g�섎���M���飾�z��>�g�rR5��1��7۽P   P   XMŽ௢�*�G���]���Gˍ������^Ž�3���� ���O�Ž���8��N���M���7��'���ӏO��� �� ��P   P   ��׽sl��1\��O����T���Za��xq����׽>	��/��H_��k���8����<��*q���Q_���/�o	�P   P   �5�8����1���&��A��������&��O/��M����&�cE���5��H_�Ž��섎�q����Ƃ��]_�Ϯ5�!R�P   P   a�B���A ���錽R���
�{����[䌽*����w����cE��/���O���g�	q���g�S�O�0��Z�P   P   �N彮���&���[����ځ�h�w�Z�w��ԁ�oy��G����w���&�>	��� ��i5�k�A���A��|5��� �|+	�P   P   3 ؽwչ�.���������+�u���p��u���oy��*���M�����׽�3���F�'���������Z��`��P   P   �Ž����M��C���D䁽�u� �n���n��u��ԁ�[䌽P/��yq���^Ž[۽�������_��B۽P   P   ����ߢ�����A��������w���p���n���p�Z�w�����&��Za�������氽�ɽ�w�ƽ�Dʽ�ƽ�佽P   P   1����Õ�xꍽ�������|���w��u�+�u�h�w�
�{������Gˍ�6���5y���㣽�����������P   P   ~ ��pމ�������r���������D䁽�����ځ�R���A����T��]���y����É�
쌽E���&��	P��P   P   S'�����Q���ށ�������A��C������Z����錽�&��O���G���s����v�����'���B��H��P   P   MPn�,�q�e�w�Q������xꍽ����M��-��&���A ���1��0\��*�7���Cq����w��q�3:n�R-m�P   P   �c��Yh�,�q����pމ��Õ��ߢ�����vչ�����A���8���sl��௢�m�����������q��6h���c�P   P   ��7�o;��JG���[�ez�k���G��V�ýS�۽݄�����c���۽�9ý;���͐���y�Q�[�MG��R;�P   P   �R;�3b;��F��M\���[��������9�LD�,��T��2���x�N���߽D��m����H���[�Q�E�P   P   MG�"e@�.4G��B\��倽Y~��B[Žm������7��SN���V� 6N��~7����32����Ľ44��ӯ����[�P   P   Q�[���J���J�^�[�ң�!w����ɽ�h��l*�L�V���������~���c��TV��+*��/�Kɽ54���H�P   P   ��y��Y[�l�Q�
{[�Y�y��䘽\IŽZb�"�0��oi���������0������}���)i��K0��/���Ľm���P   P   ͐�L#r�f\��t\��Pr���h|���~���\*��di�$Z��sI¾�ܾ�ܾ�/¾�:���)i��+*�32��D��P   P   ;����[��i�j��_��j��s��+"������UzV�i���NC¾�,뾸�� ��/¾�}���TV������߽P   P   �9ý�~��K4|�e�.e�ZM|�|���\Sý"'��7�r����ܾ�������ܾ����c��~7�N�P   P   ��۽8����o��)�l�5�a��l�dx��w����۽�x��/N�2x��(��ܾ�,��ܾ�0���~��!6N��x�P   P   �c���������ݼt���`���`���t�����A����R�Ԩ���V�3x�����NC¾tI¾���������V�3��P   P   ���5�����9�{��a��<Y�	�a���{�%������j��Ԩ��/N�r�i���%Z����������SN�U��P   P   ބ� B��A������b�H�T���T���b���� ,������R��x��7�VzV��di��oi�M�V��7�-��P   P   T�۽#Ҵ�+�����c�I�R�^�M�u�R��b����%���A����۽"'����\*�#�0��l*���MD�P   P   W�ýd������R�{�|�b�k�R�|K�nwK�u�R���b���{�����w���\Sý���~��[b��h�n����9�P   P   �G��������T�t���a�i�T�5�M�|K�^�M���T�	�a���t�dx��|���+"��h|��]IŽ��ɽC[Ž����P   P   k��z����|�W�l�ma�/bY�i�T�k�R�I�R�H�T��<Y���`��l�[M|��s���󐽆䘽"w��Y~��\���P   P   fz�R�r�k�&]e�:b�ma���a�{�b��c���b��a���`�5�a�.e��j��Pr�Z�y�ӣ��倽��P   P   ��[�D�[���\�(�_�%]e�W�l�T�t�R�{�����8�{�ݼt�)�l�e��_��t\�
{[�_�[��B\��M\�P   P   �JG��K��R���\�k���|��������*��A����������o��K4|�h�j�f\�l�Q���J�.4G��F�P   P   o;���@��K�C�[�Q�r�y�������d���#Ҵ�B��5������8����~���[��L#r��Y[���J�#e@�3b;�P   P   �����������/��8R���������\�����ݽu�������/d���fݽ�@������X���Q�TR/�������P   P   ������8{�I0���X�]#�����H㽚���h#��v1�f1�M<#����H�����Dʉ�t]X���/��E�P   P   ���x=�����=0�bX[�#���	���]i�d�)��WS��t������Zt�3S��6)� ��V��xB����Z���/�P   P   TR/��������/�"�X�,����7ƽN�
��i@�j{���Q��`������l(��I��@���
���ŽxB��t]X�P   P   �Q�y�.��2$��!/�OR����C���Y�
�I�莾�������� ��s���������H���
��V��Dʉ�P   P   �X��?I�l0�-0�Y<I�:����IT��S@��ߎ�j*ξg�
�n�$�4�$�}�
�:�;����@� ����P   P   ���I�j���@���3�W�@���j��Ν�;��bd)��f��#���ʢ
�5�`�H���4�}�
����I���6)�H��P   P   �@��f����]U�'�:���:�1U�����d�����0'S�6��G��x�$���H�`�H�4�$��s�m(��3S����P   P   �fݽ�3��5�k�nD���7��)D���k��B���sݽ�>#��Tt� �� �x�$�5�n�$�� ������Zt�N<#�P   P   0d��d����I��GaN�N�7���7�iN�=M��?����R���Q1������G��ʢ
�g�
����a������f1�P   P   �������J����EW��9��m0�֠9��AW����ﵽC����Q1��Tt�6��$���k*ξ�����Q���t��v1�P   P   v���,��Gz���|\���;�x�,�߄,��{;��i\��e��ﵽ�R���>#�1'S��f���ߎ�莾k{���WS��h#�P   P   ��ݽ���Dχ���\�sR<���*���%���*�	B<��i\����?����sݽ���cd)��S@�I��i@�e�)����P   P   ^����o���m��{mW���;�7�*�#V#��R#���*��{;��AW�=M���B���d��<��IT�Z�
�O�
�^i�I�P   P   ����ވ��(l�m�N���9�@�,�l�%�#V#���%�߄,�֠9�iN���k�����Ν��D����7ƽ
������P   P   ����k�:�U��aD��8�9�0�@�,�7�*���*�x�,��m0���7��)D�2U���j�:������-���#���^#��P   P   �8R��uI��A�G	;�� 8��8���9���;�rR<��;��9�N�7���7���:�X�@�Z<I�PR�#�X�cX[���X�P   P   ��/��S/�xl0�}04�F	;��aD�l�N�zmW���\��|\��EW�GaN�nD�'�:���3�-0��!/���/��=0�I0�P   P   ���3���s$�xl0��A�9�U��(l��m��Dχ�Fz��J����I��4�k��]U���@�l0��2$������8{�P   P   ���e�3���S/��uI�k�ވ��o�� ���+�����d����3��e���H�j�?I�y�.����x=����P   P   2塼�x����ż�$����!�9ZW�ݍ�aᴽ��ڽ0S���� �����ڽ�u���u����V�;!��Y���+ż.9��P   P   .9���]��4ü����J)�0m� ���{%�|��00�@�B��B���/����ύ�"���Gl���(�����0�¼P   P   �+ż�o����ż����,���y��@��$d��38���p��������������Zp��7���𮶽��x�4�+�����P   P   �Y��}�ͼF�ͼ�����3)���y��ν�MV�i�V������Ⱦ�n�aS�fKȾ"r���ZV�����>����x���(�P   P   ;!�Z����ݼ|����!�&�l�%)���L�C�b�T	��B���%�޲7�e�%�x�������B=b����񮶽�Gl�P   P   ��V�(�����<��3���W�9k���J�ݿV�w����	�xhM��悿Wق��.M�k|	������ZV���#��P   P   �u����=����K� ���&>�ʰ��M�ཀྵ8�r��������]M��t���Ŭ��`���.M�y���"r���7�ύ�P   P   �u��0�j��&�s	�&$	�0�&���j�����ͧ�@�p��dȾJ�%��Ⴟ�ɬ��Ŭ�Xق�f�%�fKȾ�Zp����P   P   �ڽd���@�e��Y>�~��A��y��_�ڽ �/�����I�c�7��Ⴟ�t���悿߲7�bS�������/�P   P   ���/����cY��S!� ������a!�TrY�����u����B�i☾�I�J�%��]M�yhM��%��n������B�P   P   �� ��[���k�^I,�G��<�>�JK,��k�VE���� ���B�����dȾ�����	�C����Ⱦ ���A�B�P   P   2S��/m���q���2�q;����������8�o�2��wq�VE��u�� �/�A�p�s���x���U	��	�����p�00�P   P   ��ڽ0'��O@k��2��|�
:��a?�4��ts�o�2��k�����_�ڽͧ��8�޿V�E�b�k�V��38�}��P   P   bᴽc����Y�@p,�L��D����%�4���8�JK,�UrY��y������N���J��L�NV�%d�}%�P   P   ݍ�*k�BA�ڍ!��9�i���J���a?�����>��a!�A���j�ʰ��:k��&)���ν��@��!���P   P   :ZW��G>�'��������V�i���D��	:�������<������0�&�'>��W�'�l���y���y�2m�P   P   ��!���-8��]	�Sr�����9�L��|�p;�F� ��Y>�&$	���4���!��3)��,��J)�P   P   �$�����N����� ��]	����ڍ!�?p,��2���2�^I,��S!�e��s	�K� ��<��}�������������P   P   ��ż�
μ�G޼N���,8�'�BA��Y�N@k��q��k��cY��@��&��������ݼG�ͼ��ż5üP   P   �x�������
μ������G>�*k�b���/'��.m���[��.���d��/�j��=�(��Z��~�ͼ�o���]��P   P   G���!�»���k����Ѽ+p#���o�$I��"\н���Y����K�Ͻ�ϣ�6�n�J�"���м�~�^������P   P   �����Q»��Xʁ�D���;��V���׽.�y�7��N�8�N�S�7�X���iֽ<��#:���Y�����P   P   ^�����
���������EI�h�����A�A�G���u<���x���W��X7A�Ri�����H�.��Y���P   P   �~���(�T)���������H��쭽W�@ h�OR����.N��8����ꮾZxg�С��D��H���P   P   ��мQ�|��RK�T�}��Ѽ��:�O��=��<w��̾�� ��oc�RT��U+c��E �Y̾ʔv�С������#:�P   P   K�"��޼� 1��a��r���6#�`.��^����g�w̾�3��v���̿2�̿&?��ݧ2�Y̾Zxg�Ri�=�P   P   7�n�_5��۫��ލ�U.�����,_o���ֽ4�A��-��� �Tn������������&?���E ��ꮾY7A��iֽP   P   �ϣ��5:�P/ἐx��󙢼܏Ἔ�:�0��_���t�����Nc���̿����3�̿V+c�­�W��X��P   P   L�Ͻ�Zn��H�by���l��0���6s�ȓn��нn�7�����5�CO����̿������̿ST���8�y��T�7�P   P   ��a~��s1*�_ݼ������>ݼ_H*�4���]��2�N�^����5��Nc�Un���v���oc�/N�𞯾9�N�P   P   �Y�� ���wj>�f���������<!��>����g>�N����$��3�N�������� ��3��� ���w<��	�N�P   P   ���L����E�Bk������1���7��U���f�0�E�O���]��o�7��t���-��w̾�̾QR��H���z�7�P   P   $\н����n�>��x�)D¼�ӟ��o���ן��B¼f��g>�4����н`��5�A���g� =w�A h�C�A�/�P   P   &I����n��*���������@ן����Ò��ן�U���?���_H*�ɓn�1����ֽ_��>�Y�����׽P   P   ��o�u�:�ͨ�K~ݼ@A���B���p�����o���7��<!���>ݼ6s���:�-_o�a.��O���쭽h���V��P   P   ,p#����<��o�3���.��B��?ן��ӟ��1���������1���܏Ἂ���6#���:���H�GI��;�P   P   ��Ѽ�ν�m������O���3��?A��󥾼(D¼�������򩼑l��󙢼U.��r���Ѽ������F��P   P   l��J~��Ƃ��S�����m�I~ݼ�����x�Ak�d���^ݼay���x���ލ�a��U�}��������Yʁ�P   P   �����)��5L��Ƃ�l���:��̨��*�l�>�
�E�uj>�q1*��H�O/ἅ۫� 1���RK�T)�����P   P   "�»��ﻢ�)�J~��ν����s�:���n�����K������`~���Zn��5:�_5��޼�P�|���(�����Q»P   P   ��5<�C$<�E�;T��9�L#��\̼��7��ŋ�����}��q����.����E����6���ʼ�!���9�)�;%�$<P   P   &�$<'m$<b�;�8g�B�s~��Oo�Kk½M���6��P�2�P�E6���������m�����- @�0ec9���;P   P   �)�;�P<.��;�� 9��N�����ow��[|A����7E���&�����̴����@��}���8�����L�(ec9P   P   ���9y
�;�B�;ș9mB����,���
��zm��Ƽ�ܧ�~�'��'�h�G��εl�3
�N����. @�P   P   �!�;��9��`;���9��"�~1��֌��
�  ��k��<��ǋ��T�������=<���߾�8~�3
��8������P   P   ��ʼ�0��A#��]��������˼^�n��;���Tm�{Y�`�U�-W�����r������)U���߾ϵl��}����m�P   P   ��6��������������d@��>57�$½{CA�������<��K���4�i�e��c4�����=<�G����@����P   P   �E���� ��aT�����Z6���8U��%�I�������ى�����������E�e�i�e�r������h�ʹ�����P   P   /����%9��d������4Ļr��˫�:j9�5����V6����i�'�hS�������4� ���T���'����E6�P   P   ��c�i�F���b� ����(��ob�C���i����V�P�<
��j�'������K��.W���ǋ���'��&��4�P�P   P   s��� ���
����Խ�.,�����A7��g�
�R��"��V�P���������<�b�U��<�ݧ�8E���P�P   P   ���4�����O"��s;���E���+;�.�����R�� ��V6��ى�����|Y��k��Ƽ�����6�P   P   ����kj�$�
�D8���E�),	��U�iK	���E�.��g�
���i�5������|CA��Tm�" ��zm�]|A�O��P   P   �ŋ�ڻ9��t�PK��t;�o*	�vk�)��iK	��+;�B7��D�:j9�J���$½�;���
��
�rw��Mk½P   P   ��7��f���R�b�H�����%�uk��U�E�����ob�˫��%�?57�`�n�֌�-���Ro�P   P   �\̼����̽U��H�7j��I)����n*	�(,	���-,���(��s���8U�f@����˼�1��������w~��P   P   �L#�e����»���?�Ļ5j��F��q;���E�p;�ҽ�����4Ļ[6����������"�mB���N�k�B�P   P   ��9�!�9��ƹ�������H�N�b�NK��B8��M"������b����������w���{��9/̦9� 9��8P   P   �E�;R�;E�];p�ƹ�»ȽU����t�"�
�����
�C�輤d���aT�����4#����`;�B�;+��;_�;P   P   �C$<.�<R�;�!�9]���񘗼�f�ػ9�hj��4��� ��a�i��%9��� ������0��K��9y
�;�P<&m$<P   P    ��<��<��<�<H�;JV
�X0켁�Y�U����Ž�"Խ`JŽ����;�X��h�؂���;��<[�<d��<P   P   d��<A��<*��<�Y�<���;��e���,�7���uG��wE+�<�F�[�F���*��x���;����+�7b�K��;j�<��<P   P   [�<H��<��<�]�<Bc�;�鎼f�W�Ebؽb=6�����Ь�q���З���8���5��d׽�{V�,���<d�;i�<P   P   ��<f��<Oʴ<��<��;3ӎ��?h�����Md�t����	�YK,�5*,��	�剻���c�� ��X�f�-���J��;P   P   ��;b��<�_�<!�<�o�;�Ne���W�% ����v����K�B��&���⪿�푿�EB�6(�,�u�� ���{V�7b�P   P   ڂ���<�+�<H�<��<s�	��,��&ؽ&d����r]�m4̿��������˿��\�6(ᾗ�c��d׽��+�P   P   �h�^�"�,d<�W<ۨ<��(�#������6�廾��B�*̿hbC� �y�#C���˿�EB�剻��5��;��P   P   =�X������;J3<!�<���:�j���Y�,���_���	�������Sz�!�y�����푿�	��8���x��P   P   ��8e��Zػ�i�;E��;[{�;ڻ���������+�����/,��窿���hbC�����⪿6*,�З����*�P   P   aJŽ��/�F�p�V,f�i��;ɢ�;��m��jq���/��CŽ��F��q���/,����	*̿n4̿�&��ZK,�r���\�F�P   P   �"ԽB�M��|�����U��:ғm;e��:U�������RhM� �ӽ��F�����	���B�r]�L�B���	��Ь�=�F�P   P   �Žq�M��/��O� �g�(��;;�;H�-����"��ShM��CŽ�+��_��廾��ᾉ��u�����yE+�P   P   W���B�/�=Ũ��� �~}ź��:��:��:�:Ⱥ��������/�����-����6�&d���v��Md�c=6�wG��P   P   ��Y�{��X�q��4���'����:<�:��:��:L�-�W����jq������Y�����&ؽ' �����Gbؽ9���P   P   ]0��Ƅ���ڻ�k�>p�:�,;q�:@�:��:�;b��:�m�	ڻ�j��%���,���W��?h�i�W���,�P   P   PV
���*���:<��;k$�;��n;�,;덜:
�:�;;ԓm;ɢ�;Y{�;���: �(�w�	��Ne�6ӎ��鎼��e�P   P   ?�;s<D�<��<7��;m$�;Qp�:ą'�f}ź>�(�e��:k��;E��;!�<ڨ<��<�o�;��;:c�;���;P   P   �<\�<9�<�xW<�<B��;��k�{4���� �J� ����),f��i�;K3<�W<G�<!�<��<�]�<�Y�<P   P   ��<	��<�*�<:�<F�<8��:��ڻQ�q�9Ũ��/���|��A�p�Zػ�;-d<�+�<�_�<Nʴ<��<)��<P   P   ��<	��<	��<]�<s<��*��Ƅ��z��?�/�n�M�?�M���/�5e������T�"���<b��<f��<H��<A��<P   P   ��1=�-=�I!=[�=���<ڮ<�XK��M���y����ᵽ}���i7~�j�B4H��	<�q�<�$	=�o!=E�-=P   P   E�-=-�-=%�"=�u	=V�<�X;�Dͼ�����޽C���c7�E7�CK�� ޽p[��˼`�e;⋶<f�	=�#=P   P   �o!=Si(=�I!=�r	=��<g�79�8�����%��z|�
�����������b�{�-K%�e!�����m�9
(�<f�	=P   P   �$	=�=�=��=���<��@9�1 ���ֽ&�S�J��|w��!�-� ��;��ѱ���R�X�ս��m�9⋶<P   P   �q�<�0=n=X�=_��<�Z;�� �ֽ��e�?E־�4�����bu���`���^4��վ�"e�X�ս���[�e;P   P   �	<���<u!�<���<� �< �<�̼�ϵ�I~S�a2־BL�_ϱ�� �h����y��&�K��վ��R�f!��˼P   P   E4H���U<�V�<��<W��<'DT<)}J�Ɂ�2�%�X��u�4��Ǳ��T��fF��"��y���^4��ѱ�.K%�q[��P   P   j���e��<�W�<3�<�2�<7'�����&n޽�|��V�T��� ��yF��fF�i����`���;�c�{�� ޽P   P   k7~�z�6|�;"��<�^�<NF�<���;�r��mp~�PQ������� ��x��� ��T�� �bu��.� �����DK�P   P   ~����\�ۼ	�<]&<�oq</:q<0�%<KO�b�뼉����!7�xв��� �U���Ǳ�`ϱ������!�����E7�P   P   �ᵽ3��
����;%+<�[B<��*<T��;k
�l��$����!7������V�v�4�BL��4�|w�����c7�P   P   {������G0�n��:`��;��<�<���;�D�:�W0�l������QQ� |�Y��b2־@E־J���z|�D��P   P   ��'�;~
�_��:!�;���;l�;D�;E��;�D�: k
�c��np~�'n޽3�%�J~S���e�'�S��%���޽P   P   �M��ق��M�U��;0�;��;ϟ�;F9�;D�;���;R��;UO��r�����Ɂ��ϵ�"�ֽ��ֽ������P   P   �XK��4����;|e&<�s+<�e<���;П�;m�;�<��*</�%<���;V'��.}J� �̼���1 ��8��DͼP   P   Ӯ<:8T<�W�<z��<G�q<�	C<�e<��;���;��<�[B<.:q<MF�<�2�<$DT<��<�Z;a�@9Ζ79�X;P   P   ���<\�<^%�<�m�<S��<I�q<�s+<6�;'�;e��;'+<�oq<�^�<3�<V��<� �<]��<��<��<T�<P   P   [�=o=��<k0�<�m�<{��<�e&<_��;���:���:���;>]&<#��<�W�<��<���<X�=��=�r	=�u	=P   P   �I!=��=�=��<_%�<�W�<��;M�4~
��G0�
�ȼ	�<|�;f��<�V�<t!�<m=�=�I!=%�"=P   P   �-=�_(=��=p=]�<@8T<m4���ق�!�
��0���\�w��􀺘�U<���<�0=�=Si(=-�-=P   P   m=��i=��]=rhF=��=���<*[�:�"Ƽn�O�B����"z����N�O�ļ�f ;ԕ�<]=7�F=��]=��i=P   P   ��i=b�i=��_=��H=&�=u�<D$��#N�ɽk�M0��10�e���gȽ�L��m ��`�<�=v�H=��_=P   P   ��]=!�c=	�]=�xH=�J=~��<�.�����u���w��ʡ����F�v��a��N���ޠ��;�<��=v�H=P   P   7�F=$+W=XW=-SF=�=�Æ<o�¼�ʽ��IL��+��@? �@7��#�. ��˯�S�K��켽�{���;�<�=P   P   ]=��@=��I=�j@=5�=�$�<{Ԣ�����O_���Ӿ�,���q�����n�q���,��5Ӿc|^��켽�ޠ��`�<P   P   ԕ�<�>=�k4=V4=��=ګ�<�@#��֛��L���Ӿ;@����M�˿D�˿�嚿�?��5ӾS�K��N���m �P   P   �f ;_�<��=�� =��=z{�<:'�:T�M�<��>����,�p	���������f�嚿��,��˯��a��L�P   P   R�ļ�4=< ��<�=�={�<<<T?żφȽH�v�E �Y�q�N�˿������E�˿o�q�. �G�v��gȽP   P   ��N���T��</��<���<A��<�-�<�f���N���y����
�r���N�˿���M�˿�����#��f��P   P   #z��烓�L��;xg�<fB�<�%�<�"�<zg�;}���F��)�/�gٰ��
�Y�q�p	�������q�@7����10�P   P   ������ռ�(����0<��j<G�u<�1j<�0<�����pռ&��*�/�y���E ��,�;@��,�A? ��ʡ� M0�P   P   D����ּ��-���;H�#<�(<��'<d#<��;D.��pռ�F����I�v�?�����Ӿ��Ӿ�+���w�l�P   P   q�O����JV���I�;�1
<C��;��;���;di	<��;~���
}���N�ІȽ<���L�P_��IL�v��ɽP   P   �"Ƽ�����;?�0< $<�z�;&��;�e�;���;c#<�0<sg�;�f��W?żV�M��֛������ʽ�����#N�P   P   �Z�:v�;<v�<��<^gk<-�(<���;'��;��;��'<�1j<�"�<�-�<z<<'�:�@#�Ԣ�s�¼�.��D$�P   P   ���<U��<P��<�J�<ʧ<}�v<-�(<�z�;E��;�(<G�u<�%�<@��<{�<x{�<ث�<�$�<�Æ<|��<s�<P   P   ��=�!=x�=>�=hR�<ʧ<agk<$<�1
<K�#<�j<fB�<���<�=�=��=4�=�=�J=%�=P   P   qhF=�@=ڄ4=w� =?�=�J�<��<D�0<�I�;��;��0<yg�</��<�=�� =~V4=�j@=-SF=�xH=��H=P   P   ��]=�.W=
J=ۄ4=x�=R��<v�<�;�R����-��%��T��;U��< ��<��=�k4=��I=XW=	�]=��_=P   P   ��i=&�c=�.W=�@=�!=X��<}�;<o�������ּ��ռ䃓�	���4=<`�<�>=��@=#+W=!�c=a�i=P   P   K�=�|�=E�=M�x=�O=>�=�.5<������D����v
��'����dD�����u7<J�=3=O=Ӛx=�=y�=P   P   y�=lw�=�F�=�}=��P=z� =,𔹴#;���νJ���@���@�:
�QXν7:����A_=�6Q=�'}==L�=P   P   �=�W�=Uڇ=��|=$�P=);�<�}*�;���O�(��]���s����ʾgM���#���h(��ٗ���&��t�<ARQ=�'}=P   P   Ӛx="Q�=4J�=_nx=%�P=1D�<��l�վ���`���ɾ�;z6�fk6�����Mɾzp`����q�h��t�<�6Q=P   P   3=O=V�m=��u=]�m=��N=� =U�)�����Qw�E���YJ�����㌜��勿�/J�����v������&�A_=P   P   J�=>XG=D [=��Z=�#G=�y=�a��3����`�P!����`�R�����߿,�߿D���(�`����{p`��ٗ�E��P   P   t7<85=��5=a�>=r�5=��=��5<�Y:�gq(�Gɾ�#J����fN��z���O��D����/J��Mɾ�h(�7:�P   P   ����Bw�<��=��=9�=q�=��<�摼�1ν� �� ���ǋ���߿���z��,�߿�勿����#��RXνP   P   �dD��1�:���<;<�<}��<��<y�< Y�:LD���� ����6��\����߿fN����߿䌜�gk6�hM��:
�P   P   (����>j�hV<^��<n�<(�<�W�<��<��i�����X@�Nsʾ�6��ǋ����S�������;z6���ʾ��@�P   P   w
������
�:�o<�O*<��%<��)<��<�n�:�ҿ�Ls���X@� ��� ���#J���`��YJ���s����@�P   P    ���߼����ͺz-�;��;�94;�3;��;��;��ͺ�ҿ�������� ��GɾQ!��E����ɾ�]��J�P   P   ��D��k��Ȼ:���;�a;T絺 C������\;��;�n�:��i�MD��1νgq(���`�Qw���`�P�(���νP   P   ����)��:ʒ<�<zd�;늲�a㥻��������}��;��<��<�X�:�摼�Y:��3������վ�<����#;�P   P   �.5<=0�<\��<�#�<��+<c�8;X@�a㥻 C��3;~�)<�W�<y�<��<��5<|�a�[�)���l��}*��P   P   =�= .=�+=���<���<�'<f�8;⊲�M絺�94;��%<'�<��<p�=��=�y=� =/D�<';�<y� =P   P   �O=PiG=z%6=h6=���<���<��+<d�;�a;��;�O*<n�<|��<8�=q�5=�#G=��N=%�P=#�P=��P=P   P   M�x=�n=?G[=��>=h6=���<�#�<<��;�-�;�o<^��<;<�<��=`�>=��Z=]�m=^nx=��|=�}=P   P   E�=c�=��u=?G[=z%6=�+=^��<В<�Ȼ:��ͺ/�:kV<���<��=��5=C [=��u=3J�=Uڇ=�F�=P   P   �|�=d�=c�=�n=QiG=!.=@0�<g��:�k�ۼ�������>j��1�:Bw�<85=>XG=V�m="Q�=�W�=lw�=P   P   �D�=���=��=��=cNm=r#=iZY<�ݫ���k�Ռ��ÄȽ*]��5k�(ݪ�`�Z<P�#=~:m=�Ռ=��=���=P   P   ���=<��=c��=��=��t=�=y�;@|V��<��v�C��~q��cq��VC����#vU�;xb=�u=���=���=P   P   ��=]Ӛ=��=$ِ=��v={==JI��/���P��R��3�tk�q��6��(P�u~����	�1�=Mw=���=P   P   �Ռ=!y�=wu�=�Ɍ=��t=|?=^�V�!��`����q��bN�+�����;N�"H�Gt�����/pS�1�=�u=P   P   ~:m=*�=�=���=�m=�=�2�sὩ朾�.%�S����ο���>	ο�w��%���������	�yb=P   P   P�#=�H[=�j=��j=�%[=�P#=�;[���~��x%��>�����h�(�a�(����A��%�Gt��u~��;P   P   `�Z<f{=m�;=��A=��;=eZ=xZ<OeU�;P�*��W������?�)�Y��?����w��"H�(P�#vU�P   P   )ݪ�5C�<��=�=Â=Zj=�'�<�q��%������/�M�d�Ϳ��(�H�Y�)�Y�a�(�>	ο�;N�7�����P   P   5k����p�<L!�<��<���<WR�<@�/lj���B�IL񾘸��NY迚�(��?�i�(������q���VC�P   P   +]���K����:;_��;���;�\�;�;��:;Az�������p��������d�Ϳ�������ο+��tk��cq�P   P   ĄȽl��m~�55��A��o�ѻ���^P7�V��� ���ǽ�p�IL�/�M��W���>��S����bN�3�~q�P   P   ֌��Ւ�< 1��)��&Z� ���+����Z�z���0�� �������B�����*�x%��.%��q��R��v�C�P   P   ��k�������l��wX���$����ؼ0�������{��[��Cz��0lj�%��<P�~���朾`����P��<��P   P   �ݫ�����=;��0��+Y�5����z�F��0�����Z�jP7���:;.@��q��QeU�[���s�"�Ὦ/��A|V�P   P   dZY<�U�<��<7<=|���=���pؼ�z��ؼ�+������;UR�<�'�<rZ<�;�2�c�V�OI�d�;P   P   r#=ު=�=9I�<$��;%�̻�=��4����$�� ��s�ѻ�\�;���<Yj=cZ=�P#=�={?=z==�=P   P   bNm=N�[=KC<=.=py�<'��;8|���+Y�vX���&Z��A�����;��<��=��;=�%[=�m=��t=��v=��t=P   P   ��=�-�=nk=�iB=.=;I�<7<t�0�h���)�55�^��;K!�<�=��A=��j=���=�Ɍ=$ِ=��=P   P   ��=���=|%�=nk=LC<=�=��<��=;���7 1�f~껨�:;�p�<��=l�;=�j=�=wu�=��=c��=P   P   ���=��=���=�-�=O�[=ߪ=�U�<�����Ӓ�j���K��
��5C�<e{=�H[=*�=!y�=]Ӛ=<��=P   P   �˧=��=�̟=�a�=�r=�)=�*�;1
�3c��\�����'�4����	���;�= dr=3�=֣�=���=P   P   ���=���=�â=O�=�z�=$�"=N-�f���,� �&*~����Z���}�� �����w�$� �"=�m�=�֘=گ�=P   P   ֣�=��=��=��=sу=Z�=�,e��B����W�&�I.:���%����φ���ub��; =Ӄ=�֘=P   P   3�=�M�=]N�=(4�=�c�=��=#Қ��R��乾M�8�$	���*�����J쓿�m8��������.e���; =�m�=P   P   dr=B�=W�=[@�=mSr=_�"=��c��.��Ͼm�h��ֿ@[�{�1�R���տ�eh���ξ���ub� �"=P   P   �=�Q=s�\=��\=1�Q=#�=|�&������^h�W����I�$��.����I����eh�������r�$�P   P   ��;A�=�=�� =�=�=���;�ǌ�ߧ���78���տ\�I�S<��蛩��J����I���տ�m8��φ�����P   P   ��	� 7<���<���<��<J��<�<SM	�# �	z뾨��������1���蛩�.��R�J쓿��� �P   P   4������7;�:8%;�>�:��$;�%�:����|����|�	n%������>1����S<��$��{�1������%���}�P   P   �'�6�F���}����U*��6 ~� ���Wq�~��O���~9�������\�I���I�@[��*��I.:�Z�P   P   ���p�U���H,�����Q ����)d��D�s�T�i!��O��	n%�������տW���ֿ$	��&����P   P   \�E�U��
�����LD��b���b���D����b�	�t�T�~���|�	z뾗78�^h�m�h�M�8�W�&*~�P   P   4c�����7�V���WU�'����7���Ƀ���U�����D�Yq��|��$ �৆�����Ͼ�乾���,� �P   P   1
������]���Q�s�C����V��c1���Ƀ���D�*d�������UM	��ǌ����.��R��B�g���P   P   �*�;�*<9\�:n{�� ��Qb����V���7����b����; ~�O%�:�<���;��&���c�$Қ��,e�N-�P   P   �)=�a=A�<c�2;e������Qb����'����b��Q �W*����$;F��<�="�=]�"=��=Y�=#�"=P   P   �r=mgR=<�=쌲<�~�:e��� �r�C��WU��LD��������>�:��<�=0�Q=lSr=�c�=rу=�z�=P   P   �a�=��=N]=�!=팲<n�2;j{��Q�U����G,��}�8%;���<�� =��\=Z@�='4�= ��=N�=P   P   �̟=��=�`�=N]=<�=C�<a\�:�]���7��
���F��+;�:���<�=r�\=V�=]N�=��=�â=P   P   ��=�-�=��= ��=ngR=�a=�*<�����D�U�o�U�5�����7<@�=�Q=B�=�M�=��=���=P   P   ��=ϡ=�;�=FZ�=�xZ=Z��<�ܻ�ha��޽�s��..��W�;A޽z'a�e4ݻ���<��Y=��=���=���=P   P   ���=��=;��=���=olw=��=u�[������I�«��T�žΧž�{��ueI������<Z�؂=4w=�m�=`{�=P   P   ���=-ܚ=��=G��=%'�=��=>v¼�$�.t��U��p���T�8;�t���~��R����=B�=�m�=P   P   ��=�_�=oe�=Y�=N,w=��=����/��S羻�m�1�ÿw���iy��	�ÿ?m���R'/�Љ輓�=4w=P   P   ��Y=�i=�Tj=#�i=��Y=�~=���1b/�k��sy���X��eS��q�{VS�D��X��;`�R'/�Q��؂=P   P   ���<�$=�(=[$(=� $=��<;Z�������W��A�"�~i���а�Ѱ�
j��b�"��X����~���<Z�P   P   a4ݻu�<���<�ע<���<WD�<3Oۻe����c����l��"�T��h��lz���+��
j��D�?m�s�������P   P   y'a��
9�L�w�j����-v�|8��k`���H���<ÿ�S�#���5r��lz��Ѱ�{VS�	�ÿ8;�ueI�P   P   ;A޽��,����I������hs�7,�Suݽp��1T�����\�p�#���h���а��q�hy����T��{��P   P   �W�������T�ޥh����f����h��]T��"��0��&�ľA'o������S�T��~i���eS�v����p�ΧžP   P   �..��_��Q���qG���U�������`���P���h��Xί��b-�&�ľ�1T�<ÿ�"�A�"��X�1�ÿ�U�S�žP   P   �s�u]��͒��W>���׽�i�9v�ؽ�X���~��Xί�0��p�����l��W��sy����m�t�«��P   P   �޽�����b���$��[�Sv������uF佀X���h���"��Tuݽ��H��c�����j���S�.�I�P   P   �ha�rh,�T�������׽�g���������ؽ�P���]T��7,��k`�f�����1b/���/��$�����P   P   �ܻ
7���׷g�c괽��w��������9v��`����h�ks�8�AOۻAZ������?v¼w�[�P   P   X��<qx�<�f��a�t���
�����g�Sv��i�����g����Lv�SD�<��<�~=��=��=��=P   P   �xZ=_�$=8Ҩ<�1��p�s���c괽��׽Z��׽�U�����	��+�����<� $=��Y=M,w=%'�=nlw=P   P   EZ�=�Xj=�-)=�+�<�1���a�ַg������$��V>��qG��ޥh�J��u���ע<Z$(="�i=X�=G��=���=P   P   �;�=��=�?k=�-)=9Ҩ<�f����T��b��̒��Q�����T����[�w����<�(=�Tj=oe�=��=;��=P   P   ϡ=��=��=�Xj=`�$=tx�<

7�ph,�����t]���_��������,��
9�s�<�$=�i=�_�=,ܚ=��=P   P   ���=�А=��=�f==n =� ><��_E�� ���E�V�Y�<�E����D������!;<�{=�'e=Љ�=g��=P   P   g��=ⵐ=7M�=���=@�O=�/�<����-�3k��浾o�R⾔����j���CU�:V�<O=�.�=U�=P   P   Љ�=���=G��=Pf�=�^=)��<*[��>!����`�(��nq�lb��u9q�[F(�%���`� ����zM�<�,^=�.�=P   P   �'e=]�e=�e=(ne=�VO=���<����C����O����߿�����&w߿ ��)� �mC���{M�<O=P   P   �{=��%=�l#=n&=o�=:��<'���C�.��(��vN$���s��Ί��xs��1$���2X�mC����;V�<P   P   �!;<��<
�<*.�<�K�<�&<<����� �
� �S���;�w�����������c�����:���(� �`� �AU�P   P   ���|R,�	9��=X�E�8�$R+��G�xn������$�L���\���5���c��c����1$� ��$�����P   P   �D����9�+�3��"H�;H��3��{9��Ϫ�uj�c�'�߿#s�����-���5�������xs�&w߿ZF(��j�P   P   �������������������ޚ��Lƨ�������!|p�wK�������\�������Ί����u9q�����P   P   <�E�3��gܽ_����f�|f�����;@ܽew�k�D���AᇿwK�#s�L���w�����s���lb��Q�P   P   V�Y���	�����d�rc-�5�5��g-��e�����	���X���!|p�߿$�;�vN$���߿�nq�o�P   P   ��E���	������'�SjF�,Y��1Y��xF���'�*����	�l�D����c�'�����S���(���O��_�(��浾P   P    ����3��;�'��:O���l�aw��l�zYO���'���ew��uj�xn��
� �.�������3k�P   P   `E���ʨ�u�۽�0��DF�ňl����.���l��xF��e�<@ܽMƨ��Ϫ��G��� ���C���C��>!��-�P   P   
��9��(�� ��w-���X�kAw����aw��1Y��g-�����ޚ���{9�����(���+[����P   P   � ><�(��P2�#A���	��l5���X�ňl���l�,Y�5�5�}f�����3�,R+��&<<7��<���<'��<�/�<P   P   <n =�z�<�2��}F��ȹ��	�w-��DF��:O�SjF�rc-��f�����=H�M�8��K�<m�=�VO=
�^=@�O=P   P   �f=�'=��<Z(R��}F�"A�� ���0�;�'���'��d�_�������"H��=X�&.�<m&='ne=Pf�=���=P   P   ��=v�f=��$=��<
�2��P2��(��t�۽3��������gܽ����,�3�9�	
�<�l#=�e=F��=6M�=P   P   �А=�F�=w�f=�'=�z�<�(�9��ʨ������	���	�3�������9�R,���<��%=\�e=���=ⵐ=P   P   �_n=�f=��J=v
=[�<
ƃ���|��!����;�g�p�^���	�p���;�;W��~�}��8��O3�<��=x�I=��e=P   P   ��e=p�e=�*]=�C=��	=���;y~C�D~�Z~�����x$�N�8|����}��V�&�C����;?�=�C=�\=P   P   x�I=�,J=�BJ=g�C={/!=��c<��;�ې(�(���@�&��sm����(>m�g]&��.��s;(��;��a<�l =�C=P   P   ��=��=�=�;=�f	=�\c<�;?�D�D�>R������e3ٿ2��y���ؿ�V�����>,D�?��a<?�=P   P   Q3�<��j<-KQ<��k<"�<u��;��;�1^D��u�����0�&l�L����l����f��#F�>,D��;����;P   P   �8��}�t����ٚ��|s��?��>aC��-(������v��V!5���x3���1��G���5��f�����s;(�%�C�P   P   ~�}��;U�Qo��w~���n�z�T��4}�y�-���o>�������0��*T���	��G�����V���.���V�P   P   ;W���@ý��ҽX������ҽf�½;����7}��	&���ؿ��k�F���M��*T���1���l���ؿg]&���}�P   P   ��;����=*�*�(�1�v*����f��p;�<ｾ�l��&��t��F��0��x3��L���y�'>m�8|��P   P   	�p�Q$7���A�xG]�Kyp�vp�4<]�ŏA� �6�b�o�a8龰y���&���k������&l�2�����N�P   P   ^���%pN�w�^�^Â��]��~���#^�����O�^�wN�@��a8��l���ؿ��V!5��0�d3ٿ�sm�w$�P   P   g�p�8eN��!i��ߍ�(饾(�����_量~卾�i�wN�b�o�<ｾ�	&�o>���v�� �������@�&�����P   P   ��;�]�6�z�^��Ӎ�|����¾*�ʾ��¾�卾O�^� �6��p;��7}�,�������u�=R��'���Z~�P   P   �!���X�	`A����OХ���¾��Ҿ��Ҿ��¾_量���ŏA��f�;���y��-(�0^D�D�D�ې(�D~�P   P   ��|�͓½�����\��/��S�����ʾ��Ҿ*�ʾ���#^��4<]���g�½�4}�?aC���;��;?���;�y~C�P   P   ƃ�l�S���ѽy�)� p�~��S�����¾��¾(��~���vp�v*��ҽ{�T��?��j��;�\c<��c<���;P   P   Y�<r�m�X�l�[��JU1� p��/��OХ�|��(饾�]��Kyp�(�1������n��|s��<�f	=z/!=��	=P   P   v
=�3q<�`��v~|�[��x�)���\�����Ӎ��ߍ�]Â�wG]�*�X�潞w~��ٚ���k<�;=f�C=�C=P   P   ��J=F=�W<�`��W�l���ѽ���`A�y�^��!i�v�^���A�=*���ҽRo� ��(KQ<�=�BJ=�*]=P   P   �f=��J=F=�3q<n�m�k�S�̓½�X�]�6�7eN�%pN�Q$7�����@ý�;U���t���j<��=�,J=p�e=P   P   g�=�=�:�<l�!<��h_�ulؽ�+�sfn�'z��𠛾~}���n�";,��7ٽ%8a�I���JR<P��<$=P   P   $=�X="=���<�<�+������!�Y���n��1-��⾳Q�������'�ሕ��𮼢><�Z�<�O=P   P   P��<�j�<���<�1�<劏<1겻Ĉp��&������h���L��e�.�L�5�G~���v&�xq��P���D�<�Z�<P   P   KR<R3�;��;�<<�<t]��ӊb�{5�Wھ�7[�m���������W����Z�C�پZG5�+�b��P���><P   P   H��������ż�կ��I��#N��yp�>\5��A�M���(S�p�@�5�[��@�L4�W`����ZG5�xq���P   P   %8a�z�x�2�����w)x�}r`��#���V&�R�پBr��o��kuz�CA���=���bz���V`��C�پ�v&�ሕ�P   P   �7ٽ��߽*����������	1߽��ؽq��QR��<�Z��(�FTz�Ok�������p���bz�L4���Z�G~���'�P   P   #;,�(�)�<��L�՗L��h<�}�'��+�󳃾r�����jL@�r%��A��������=���@��W��5�����P   P   �n��`�.2}��z��^a��/q��h
}���`�(n��ٻ��AL��	�n[�r%��Ok��BA��5�[����.�L��Q��P   P   ~}���U���]���²�an���j������%I��j.���,���q��e��	�jL@�FTz�kuz�o�@����e���P   P   𠛾p4��Ń��F�оo<꾈��o9��о�r������F���q��AL�����(�o��(S�l�����L�1-�P   P   'z��[*��h¶�&*�W��8��9��X�8-ᾫ�������,���ٻ�r��;�Z�Ar��M����7[��h��n��P   P   tfn��6��Bf����r�v��_�����{�8-��r��j.��(n�󳃾QR��R�پ�A�Vھ����Y��P   P   �+�w`��'��yVоF�P���`&��e&�����X��о%I����`��+�q���V&�>\5�{5��&��!�P   P   wlؽ��'�|�|�z��G��a"�{���`&�_���9�o9꾗���h
}�}�'���ؽ�#��yp�Ԋb�ňp����P   P    h_�aj޽?�;��#��i��R��a"�P��u���8����j��/q���h<�	1߽~r`�&N��}]��;겻�+��P   P   ���gv�
d���K����i��G��F� r�W�n<�an��^a��՗L�����x)x��I��7�<㊏<�<P   P   h�!<����h�����K��#��z��yVо��%*�E�о�²��z���L��������կ���<�1�<���<P   P   �:�<"� <����g��	d��>�;�{�|��'��Af��g¶�Ń���]��-2}�(�<�*���2���ż��;���<"=P   P   �=�j�<#� <�����gv�`j޽��'�w`��6��Z*��p4���U���`�(���߽z�x�����L3�;�j�<�X=P   P   �<��@<ѧ���U¼�k��&սY'���l��/��=���D½�ĳ��S���hm��'�hfֽ�Ln�pƼ���g�=<P   P   g�=<|�><s��;i9A�f��M]`��qٽZ&8����b���Gqؾ5lؾ����^#���g8��Lڽ�\b� J����Z����;P   P   ����1������q�G�/�,�B�������L%��g��L���!��3�!�!����zN��~b%�Ϲ�������2���Z�P   P   pƼ9�ݼ�ݼ�ļ�Ӷ��9 �e ���##�dg��m $�X\��`y���j���;����#��6��)#�������� J��P   P   �Ln�1��� LU���Om��#a��.��#�����I�F�ᵿ�F�f��	5�賵��F�Ȑ��)#�Ϲ���\b�P   P   hfֽ���2v�e�_b�
�ս��ٽ^$%�(2����F�4Ϳ�+��w_�+p_���+�!Ϳ�F��6��~b%��LڽP   P   �'��:�4�P�R�Y���P�-�:�{^'��
8������#������+�$���������+�賵���#�zN���g8�P   P   �hm��$��,X���E��=��@������Lm�����ɀﾅ�����Q_���������+p_�	5��;�����^#��P   P   �S�����������ؾ�m�b�ؾ����a���V��F����k!����A\��Q_�$��w_�f���j��!�!�����P   P   ĳ�Džq�6�50��,�Y������ľ�x����׾R3�������+��+��F�`y���3�5lؾP   P   D½��v־- �|����2��^:���2�)��J��L־-v����׾�k!��������4ͿᵿW\����!�GqؾP   P   >���f־h	�U�+���I�:a[�#a[��I��+��c	��L־�x��F���ɀﾫ�#���F�I�F�m $�K�b���P   P   �/���ľ�
���+�
DR�;�n��y���n��MR��+�J���ľV���������(2������dg���g�����P   P   ��l��e���꾹����I�H�n�����
����n��I�(�����a���Km��
8�^$%�#��##��L%�Z&8�P   P   Z'�ˁ�V���O����2��@[�.�x�����y�#a[���2�Y���������{^'���ٽ�.��e ������qٽP   P   'ս!.:��꓾rVؾ����0:��@[�G�n�:�n�:a[��^:��,�b�ؾ@��-�:�
�ս�#a��9 �E���O]`�P   P   	�k��N�rP��ӟ���ྸ����2���I�
DR���I���2�50��m�=����P�_b��Om��Ӷ�4�,�f��P   P   �U¼Y������X��ӟ�qVؾO�������+�T�+�|��5��ؾ�E��R�Y�e�LU���ļ}�G�w9A�P   P   㧎��ټ(������rP��꓾U������
�h	�, �p�����,X��3�P�1v� �ݼ����o��;P   P   ��@<Y1k��ټY���N� .:�ˁ��e���ľf־�v־Cž�����$���:����1���9�ݼ�1��{�><P   P   �,�#kn��s�R"}�ؽڈ'��ip�����PǾ6����%�ŏǾk���?4q�>X(�"�ٽ$���5�	r�P   P   	r�YUp�+��� ���o���ý���T6a�k�������גھ6�ھD
¾���V�a�Jx��HŽ%Ar���|��P   P   �5���.o�ߗ���0�����!�ѽ�.��A���Ⱦ�t��0O
��d��1Ⱦ"R���u.�w�ҽ���@�2��P   P   %������t��݌~��p�"���W���������xm� -���U�4zU���,�jB龠���B$��5�����&Ar�P   P   #�ٽى����T0���ؽ�sĽ[�ѽZ�������k���a����*Ĵ����ϰa��R����B$�x�ҽ�HŽP   P   >X(�5 ?�R
N���M���>�?�'��	��.�~��YX�%�y���ɿ?��s��V�ɿ�y��R������u.�Kx�P   P   @4q�����ǚ�E ������׊���p��<a����[龳�a�-�ɿ�>��z'�?�V�ɿϰa�jB�"R��W�a�P   P   l����ǻ���׾�j�j^� w׾�f���7k��ӽǾӻ,��埿���lt'��z'�s�������,�2Ⱦ���P   P   ƏǾӋ�4H��1��w#�%�Z1��N�,EǾ�������  U��������>�?��*Ĵ�4zU��d��E
¾P   P   �%���
�4�*��QG�SX��LX��@G��h*�ou
����.ھ(
�  U��埿,�ɿ��ɿ�����U�0O
�7�ھP   P   ��\G�/�@��k�X������{���=qk��k@�S-�C}�.ھ���ӻ,���a�%�y���a� -��t��ؒھP   P   7侷:���H��n�������Ψ��ͨ�蘙�ak����H�S-���㾌���ҽǾ[�XX��k�wm龫Ⱦ����P   P   �PǾrq
��a@�Ve������x��!AĿ�{��/��ak���k@�ou
�,EǾ7k�����~�����������A��l���P   P   ���,$��J*�Nk������n����ο��ο�{��蘙�=qk��h*��N�e����<a��.�Z������.�U6a�P   P   �ip��N����Y
G��م�	����1Ŀ��ο!AĿ�ͨ�{����@G�Z1����p��	�[�ѽ�W��"�ѽ���P   P   ۈ'�M���a׾���X��ꋿ	����n���x���Ψ�����LX�%�w׾�׊�?�'��sĽ"��������ýP   P    ؽl9>��A��#��+#��X��م������������W���SX��w#�i^辠�����>���ؽ�p���0���o�P   P   S"}�Mｖ$M�qA��#����Y
G�Nk�Ve���n���k��QG��1��j�D ���M�T0�݌~����� �P   P   �s�#~��ZZ���$M��A��`׾���J*��a@���H�.�@�3�*�3H���׾�ǚ�R
N������t��.o�+��P   P   $kn�+ �#~��M�l9>�M����N��+$�qq
��:�[G���
�ы쾻ǻ����4 ?�؉������YUp�P   P   �����$��Q��[Ͻ:� ��k��颾�Ծc7��2�����K�{e�#�Ծ~l����l�b�!���н#T��E�%�P   P   E�%�*&%��G��n����ƽ��H|M�l9��紾~پu�����VDپ�0��˘���QN�Oj�jȽː��VeI�P   P   #T����}��߀���������ɽ�t
��D�8҉�)赾�eھ�込oھ���_��!jE�w$�P"˽�3��ː��P   P   ��н�׽�׽�*нXrǽ��ɽ 꽂[�]�m��u��zc���8��N[������m�����U�P"˽jȽP   P   c�!���/��x5���/�BA!�n��"�
��\���c�L���zQ�6�f�I��6�F��ó�d����x$�Oj�P   P   ��l�셾l[��M����\"l��M���D�v�m�y����3�-mX���������`X�1��ó���m�"jE��QN�P   P   l������Ծ��۾^�Ӿ.���=#���H�����nB��2�|WX�����)3������`X�F�����`��̘��P   P   $�Ծ�	 ����N��E�J������e7Ծ-״�;�����<�5�υ��@-��)3�������6�N[�����0��P   P   |e�=9!�X.B���Z�d�K�Z��B�!�6�W�ؾ%ھ���FpI�υ����������f�I�8���oھWDپP   P   �K�Zq=�%No����ou���o������%o�7D=��\��Aa辚��<�5�|WX�-mX�6���������P   P   ���
�M�D����ѫ���ǿa^ҿ�ǿ3�������~�M�t^�\��%ھ��2��3�zQ�zc�eھw��P   P   �2���M�����Q������v�!u����G�����~�M��V�ؾ:���nB��x���L����u��*赾�پP   P   d7��>=����� B���'���W��� �|Y�;-���G������7D=�6�-״����v�m���c�]�m�9҉�紾P   P   �ԾK� ���n�w�����-N���+��+�|Y���2���%o�!�e7Ծ�H����D��\��[��D�m9��P   P   �颾�t��l�A��э�fjǿ�^��s ���+��� �!u��ǿ�����B�����=#���M�!�
� ��t
�I|M�P   P   �k�[��Lc�2{Z�Q:��$ҿ�^�-N��W��v�`^ҿ�o��J�Z�J��-���["l�n����ɽ��ɽ ��P   P   ;� ��`���pӾ�����c�Q:��fjǿ���'������ǿou��d��E�]�Ӿ��BA!�Xrǽ����ƽP   P   [Ͻ=/��ю��B۾���1{Z��э�v����A���Q���ѫ������Z��N���۾M����/��*н�����n��P   P   �Q���ֽʦ4��ю��pӾKc�k�A���n��������D���$No�W.B���Ծl[���x5��׽�߀��G�P   P   ��$���{��ֽ</��`�� [���t��J� ��>=���M�	�M�Xq=�<9!��	 �����셾��/��׽��}�*&%�P   P   ̒Z�U���0������T��Ҙ�-�о��Q�#�U>9�4A��`9��,$�hN�cyѾ�j��Y�U�U��MP��zv��P   P   zv��
1��ݿ���lƽj	��?����ݿ��|&ؾ�w���	���	�������ؾR;��֛��{�@��?
���ǽz���P   P   NP��HJ���͹�R�ƽ=�t	��0�<�f����A���rSӾ��ݾmpӾg4��V���_g���0��B
�Mw㽃�ǽP   P   V��a
����D0���	���	�ύ�L�1�϶d���c˸�U*оN1о�举F��CIe��I2�=N��B
��?
�P   P   Z�U�܃f���l�$Cf��>U��@�`60�ٙ1�s�O�����b���b�ݾU��E�ݾo���0���=P��I2���0�|�@�P   P   �j�����E����}��"嬾 ���A��3�f���d�L󇾣���? �n��F��r,�ŵ�0��DIe��_g�כ��P   P   dyѾ�V��ŷ�����X���Ѿ4֬�v������b���ﾰ��d$� ��r,�o���F�� V��S;��P   P   jN��&���@�gyP��lP�[�@���%�Q�@ؾ]ͷ�����H�ݾ�t�\$�d$�F��F�ݾ�举h4����ؾP   P   �,$��&S��;��3�����#���!��2�R�>�#��F��:Ӿ��Ͼ1���t����n��V��O1оnpӾ����P   P   �`9��z��碿%ƿ�!ܿRܿ�ƿ@Ƣ�Odz�K#9�P�	�cpݾ��ϾH�ݾ��? �c�ݾU*о��ݾ��	�P   P   4A��#������0�����������k���������A�P�	�:Ӿ�����b������b���c˸�sSӾ��	�P   P   V>9����ȿ9����7�VSU��NU���7�۳��ȿ���K#9��F��]ͷ���L�������B����w��P   P   R�#��az�N���O��	;F�S�{�����{�e<F�۳����Ndz�=�#�?ؾv�����d�s�O�жd����}&ؾP   P   ����R�D���@H��H�7�q�{�����(����{���7��k��@Ƣ�1�R�P�3֬�2�f�ؙ1�L�1�=�f�޿��P   P   .�о��%�a�����ſ����#U��ڈ���������NU����ƿ�!����%��ѾA��`60�ύ��0����P   P   �Ҙ�W���A^@�^璿��ۿN���#U�p�{�R�{�USU����Qܿ�#��Z�@�W������@���	�t	��?�P   P   ��T��s��|R���O�⨙���ۿ���G�7�;F���7����!ܿ���lP���!嬾�>U���	�=�j	�P   P   ��7}e�3J���O�^璿��ſ?H��N��8��.���$ƿ3��eyP����}��#Cf�C0�Q�ƽ�lƽP   P   �0��VL���k�|R�@^@�`���C���M���ȿ�����碿�;����@�ķ�C�����l�����͹�ܿ��P   P   U���c��VL�6}e��s��V�����%���R��az�����#���z��&S��&��V�����ڃf�`
�GJ��	1��P   P   �l��ǂ�����u�-�k��_z������̀$���H��c���m���c��H���$�?h���'������O�.�h��T��P   P   U���Ԣ�S������)�!j��0����;)����7��V �Jf �uc��i���ξgƞ��7k��*�8f��U.��P   P   j���M⽕7�wU���:�A�)��"T���������ƾ��޾��$�޾��ƾ�������U�d�*����9f��P   P   P�.�A2�)�1�6S.�A*���)� 3���I�Uo����3���AN��u]���覾Wُ��p��J���3�d�*��*�P   P   �����w���􎾪R�������}j�eJT�u�I���Q��wn�c'���d��wO��6|��5X��oo���R��J��U��7k�P   P   �'��S�Ѿ�7߾�"߾�pѾ�͹�?[��0!���Go��cn�ؠ���,������-����N��v܄�po��p����iƞ�P   P   Ah���I��'�}C-�['��������ξϠ���r���	����	:������ S���N��5X��Xُ�����ξP   P   ��$�e"M�8p�
x��xo��<	p��L��$����yzƾ����G1��X���ĕ������.���7|���覾��ƾ�i��P   P   
�H��g��l7����	ɿn�������<����H����R޾9������X���	:������xO��v]��&�޾vc�P   P   ��c��v����ֿL��z��p�q���cֿD���sc�
# �V<�9���G1�����,���d��BN����Lf �P   P   �m�������p0��\���n�Dn\��O0�����믿n{m�	# ��R޾�����	��ؠ��c'��4�����޾�V �P   P   �c�u���*�eM�P����������멎��HM�9�믿�sc���xzƾ�r���cn��wn�����ƾ�7�P   P   ��H�G������MM�^���a��X����_��f[���HM�����D����H�~���Π���Go���Q�Uo�����+���P   P   ΀$��*���Eֿ570������P��Gm��s���_��멎��O0��cֿ�<���$��ξ/!��t�I���I������;P   P   ����֥L��ि�f��/\�|r��Ӛ��Fm��W������Bn\�q�����~�L�����>[��dJT� 3��"T��0��P   P   `z�������o�X����0��|n�|r���P���a��������n��p�m���;	p����͹��}j���)�B�)�!j�P   P   k����о�&��(��$�ȿ�0��/\�����^��O����\�z�ɿwo��Z'��pѾ����@*��:��)�P   P   u�-�抾�޾s�,��(��W����f�470�MM�eM�p0�K�� ��	x��{C-��"߾�R��4S.�vU�����P   P   ��潪31�dp���޾�&���o��ि�Eֿ�����*������ֿj7��8p�'��7߾��(�1��7�S��P   P   ǂ���UὩ31�抾��о���եL��*��G��s������v���g��c"M��I�Q�Ѿ�w��@2��M��Ԣ�P   P   ��L˹��"��}E��]���4Ծ��.�>��sj���������Tх�#�j�0<?�Kq���Ծ4����mF�����l��P   P   �l�����REٽ!m�ӰA�����{k��5�����(�K6�C]6��(�va��Z�����!��f�B��&��(ڽP   P   ���� ��y�×��r!�� B�' q����_���K�ؾ��O������/پ�����'��(r���B��>"��&�P   P   �mF�ƨI�C�I���E���A�]B�~$K�b`�K1��$���'���B���(���NХ�7���{�����`�6L���B�g�B�P   P   6���jq��I���H��ޮ�������&q��`���\��&h��I|�"���&���H؇���|���h���]���`�*r��!��P   P   ��Ծi���{���c��I�ﾝ�Ծj���ɧ���)���h���c��k�Ŵt�X�t��Xl�od���h�|����'�����P   P   Mq�W�-��B�ltI���A�ĵ-��,�d�꾘w��\��� |���k��k�\�l��Lk��Xl���|�9��������Z�P   P   2<?�w�p��l������i����M��@�p�w�>�%���ؾ�\��W����lt�M�l�\�l�Y�t�I؇�PХ� 0پwa�P   P   &�j�0	���ɿ��������쿰PɿiΝ��dj�-p(��&�0���f���lt��k�ƴt�'���*�������(�P   P   Vх�(`��a��/�MjJ��ZJ���.�2��:��Ǚ��V
6������0��W�����k��k�#���D����O��E]6�P   P   ������׿f�$��o��+��Nϩ����qo��r$��e׿�ȋ�V
6��&�\�� |���c��I|�)������!K6�P   P   �����׿��0�k؎��\���2���(���C��輎�t�0��e׿Ǚ��-p(���ؾ[����h��&h�%���M�ؾ�(�P   P   �sj�;#���}$�$Ǝ� z���	y%�}�fo��輎��r$�:���dj�$��w���)����\�L1��`�����P   P   /�>�뽝����To�Y0�����@5��B5�}��C��qo�2��hΝ�u�>�b��ȧ���`�c`����7��P   P   ���Gp�ɿ�.��������i%�@5�y%��(�������.��Pɿ>�p��,�h����&q�~$K�' q�|k��P   P   �4Ծ�m-�)��A����I�������������2��Lϩ��ZJ�����M��µ-���Ծ����\B�� B�����P   P   �]���)��A��F��^o����I����X0���y���\���+��JjJ�����g�����A�G��ܮ����A��r!�ӰA�P   P   �}E�֝�����.�H��F��A���.��To�#Ǝ�i؎���o�/������jtI��c���H����E��!m�P   P   �"��H���������A�)��ɿ���}$���0�d�$�`���ɿ�l���B��{��I��A�I��y�QEٽP   P   L˹�v ��H�֝��)ﾖm-��Gp�꽝�9#���׿��׿&`��.	��u�p�U�-�f��hq��ĨI�� ����P   P   ����̽S�ބT��̞�A��b\�^�Q�H�������u훿rϔ�=*=R�Q����Mn���uU������̽P   P   ��̽fq̽]콲h�P�2�����¾A��˕��j7�g�F�+�F�١7�1������uþ�H���Q��!��=�P   P   ¡��u�hX�|���R-��P��;��([���ž(�澪/�����g���+�p�ž�롾,Ɂ�Q��!.��!�P   P   �uU��8Y��Y��U��YP�,P��FY��
n�ŗ��E����Ԩ��{����������������o��GZ��Q��Q�P   P   On���㪾���2���[��[܏��L���n�5�e�/�i���t�,���>��i��:,u�#dj���f��o�-Ɂ��H��P   P   �澖M�b�
���
�(�F澔�¾|`�����_�i�j1W�'%Q�l�P�b�P��Q��W�$dj�����롾uþP   P   S��I�>���U�{W^���U�L�>��~��L���žp���/Yt�� Q�a@�`�;���@��Q�<,u����r�ž����P   P   -=R��υ��ȟ�	�������t���?�����Q�΃��澍����T�MQP�'�;�a�;�c�P�k������+�3��P   P   ?	���k��
���Q
�M#�;���歁��97����������MQP�a@�m�P��>������g��ۡ7�P   P   tϔ�,�ܿ����S��y���x��S��L��@ܿ剔�1F�D������T�� Q�(%Q�/���{����-�F�P   P   w훿�����*E��E������3U������B���D��|��`���1F���������/Yt�j1W���t��Ԩ��/��i�F�P   P   ����^���K>U�@�� ��|����ҍ������ U��|��剔��97�~��p���_�i�0�i�F���*�澼j7�P   P   I���]Zܿ��D�^Գ����ɴ>�{�O��>���������D��@ܿ孁�̓��ž���5�e�Ɨ���ž̕�P   P   _�Q������A�����T�>���a���a��>�э�A���L�:�����Q��L��{`���n��
n�)[��A��P   P   c\��~����濥WS�2���*��i�O���a�z�O�������S�K#�>����~���¾�L���FY��;����¾P   P   A��aT>��b��v�	���x�m��)��S�>�Ǵ>�z��1U����x�P
�r���J�>�F�Z܏�,P��P�2���P   P   �̞�Q��BU�H��F����x�1���~�������������y���������U�(�Z���YP��R-�P�P   P   ބT�*E��B�
�|�]�H��v�	��WS���\Գ�>���E���S��
����xW^���
�0����U�{���h�P   P   R�@_X�\���B�
�BU��b����濐A���D�H>U��*E�����k翰ȟ���U�`�
�����Y�gX�}]�P   P   ̽��
�@_X�*E��Q��`T>��~������[Zܿ[�������)�ܿ	���υ�G�>��M��㪾�8Y��u�dq̽P   P   ;�Խ�������^��䣾7�쾱�$���Y�<���[�����rz���o���\Z��=%�������d�_�2b�C`�P   P   D`�=���5"�G[W��F����Ǿ���g"��W=�[M��%M��=���"�h��NȾ>ܓ��JX�\�"����P   P   3b�u����\"�H�3���T�)���[G����ȾCg�!%����\A�%���wɾyפ�����U�D�4�]�"�P   P   f�_��Ne�[*e�&/_���W���T��e\���p�����X��b��E��'\��|E����������q��e]���U��JX�P   P   ��:���󵾖��.0��fo�������p��@f��Gg��o�sJw���z�N�w���o��h��:g��q���@ܓ�P   P   ����� �l����U?�Q�Ǿ�F��{���C-g��O��#D��!@�wH@�B�D��AP��h����{פ��NȾP   P   �=%�kF��._��eh�A_�Z&F���$�#���ȾT0��[�n�F�C�hJ-��d&�A�-�C�D���o������wɾj�P   P   �\Z�����k��u�������?���ԋ�m�Y�jM"�(�������v���?�u<&��d&�xH@�P�w�~E��(�뾮�"�P   P   �o������������x������z���S���&���=�����ݱ�M6z���?�iJ-��!@���z�)\��^A��=�P   P   tz�������*��)h�ܴ������y�g���*�Rp�A*����L�o��ݱ���v�G�C��#D�uJw�E������%M�P   P   ������\V��C��ә��*����t��x����U�،�kĢ���L��������[�n��O��o�d��"%�^M�P   P   �[��i��Rth�{����g��F0�c=0��N��W��\"h�،�@*���=�'�T0��C-g��Gg��X��Eg뾔W=�P   P   �<������'V��y��$� ��!R���c��R��� ��W����U�Qp鿚&��iM"��Ⱦ{����@f������Ⱦ�g"�P   P   ��Y�mQ����*�E	���L�R��tv��uv��R��N�w����*��S��k�Y�"���F���p���p�[G����P   P   ��$�����G��Ӯg�JG���&0��c��tv���c�b=0��t��v�g��z���ԋ���$�O�Ǿ�����e\�)�����ǾP   P   8�쾧�E����Z��l��|j���&0�
R��!R��F0�'�����������?��X&F�S?�eo����T���T��F��P   P   �䣾�l���^�����|���l��IG���L�"� �~g�Й��ڴ��v������?_���,0����W�G�3�G[W�P   P   ��^�����$����g�����Z�Үg�C	���y��x����C���)h���r���eh�j����$/_��\"��5"�P   P   ��t�d�i��$����^����G����*��'V�Nth��\V���*������k���._�� ���Y*e����P   P   ���j��t�d������l���E�����kQ�����g������鿀������ kF����:���Ne�u�<�P   P   oN�n��;�8���m�-�����!��U�Kq�����~u��Z��T���f�U�"��i�㸥��n��39��4 �P   P   �4 �� ��,%� �6�P�^����GDþ�����C�8�DOH��bH��$9�^�����i�þ����B�_��f7�`}%�P   P   �39�?�:��8���6���=��T�;U���B����¾�������0U��=�}fþ�ʟ�3׀�^�U�o->��f7�P   P   �n��uy�5Wy�ln�F2_�&�T�8�V�E�g��`�����{٢��߫�k��������-ւ�C�h�o�W�_�U�D�_�P   P   帥�:���V*���n���o���8���^����g�k*\�qf\��Uc���j��"n�k2k���c��7]��!]�E�h�4׀�����P   P   �i�i��J��e��,����龆Yþj;��^N��LI\�X�C�ݐ7���2�Q�2��8���D��7]�.ւ��ʟ�k�þP   P   "�P�C���\���e��m\��:C���!�����ܿ¾�c��hc��g7�����:�����8���c��򓾀fþ���P   P   i�U�𳉿C��Ũ��5����٥�Xy����U��n��]�ϋ���dj�	z2���:�S�2�m2k����@�`��P   P   V����#��G���X��{�D;��?�ɷ�>U��(�8�q���es���wm�	z2������2��"n�m���3U���$9�P   P   \�����'P'�l8c�Z߆�XІ��b��'��o�6ʗ���G�F��es���dj��g7�ߐ7���j��߫����bH�P   P   �u��� ���P�W�� @��=&����������}P��| �G(����G�q���΋��hc�Y�C��Uc�|٢����GOH�P   P   ����� ��b�����2���),�I,�kg����%�a��| �6ʗ�'�8��]侲c��LI\�rf\�������E�8�P   P   Mq��[�俏�P����N[�3'M�_�M��D�����}P��o�=U���n�ڿ¾^N��l*\��`����¾��P   P   
�U�ѷ��'�鵠�vk�M�Tq�Uq�M�jg������'��ɷ���U�����i;����g�E�g��B�����P   P   �!��f��w��b�����i,��_�Sq�_�H,���� �b��?�Wy����!��Yþ�^��7�V�;U��HDþP   P   ��bC�@���������Y���h,�M�1'M��),�:&��VІ�C;��٥��:C���龈8��$�T��T����P   P   -��z��\�$B��Y/���������uk�M[�0���?��W߆��{�3����m\�*���o��D2_���=�Q�^�P   P   ��m��
��R?�Zre�$B������b�絠�}�������T��h8c��X�è����e�c���n��ln���6��6�P   P   ;�8���x����Q?��\�?���v�'���P��b���P�$P'�C��@����\�H��T*��2Wy�}�8��,%�P   P   n��̒:���x��
��z�bC��f��ѷ�Y�俛� �� ���保#���M�C�g��8����uy�=�:�� �P   P   l���B��$Y��֤��F?���߾Z���E��t��|��x��*���#Xt��)F�o��� ����튾��nP��P   P   oP��L����z�c�l���t�];��3'�������+�$9�&59��;+���ƥ����I���)wu�Km��{�P   P   ��Pч�Wt��.�l�XY�
�Y���t�y���/����Ӿ�m�r�򾠞�+�Ӿߢ��r�����u��>Z�i�Y�Lm�P   P   �튾𕾨畾Ҋ�u��Y�ߗN�*4W��o�t���G��.J�����P��~p�$X�]_O��>Z�+wu�P   P   ����л��þ/���fw��AV���u��+W�=�I��HI��>P�/�W��*[�51X���P��J�FyJ�%X���u�K���P   P   ��z[����~���8�K�߾-3�����Q|o��)I�V�2�/�'�w#�,�#�&
(��e3��J�~p�s�������P   P   !o�@^7��cO�o]X��?O�87�x������^���W�O��o'��b�|�
����&
(���P�Q��⢴�ʥ�P   P   �)F���~��D���A���1�����N~�t�E����2Ӿ����|fW��"#�Ob
�}�
�-�#�81X����.�Ӿ��P   P   'Xt�&j���ܿ������ø�M�ۿI���s���*����S���ƀZ��"#��b�w#��*[�L����꾼;+�P   P   ,���^@Ͽh��&G��Vj�J<j���F�װ�e�ο�D����8��?�R���|fW��o'�0�'�2�W�0v��)59�P   P   z�����+7����k����S��G�����#�6�(9翳Α���8���龻���W�O�W�2��>P�G���m�$9�P   P   �|��%��(E�����Fm��T@��5��7�������D�(9��D����*�2Ӿ]����)I��HI�u�����Ӿ�+�P   P   �t�O	Ͽ;�6������0�0�vPA���0��������"�6�d�ο�s�������P|o�>�I�!�o��/�����P   P   ��E��%��������ZH��N�0�fLR�JR���0��7����ְ�H��s�E�������+W�*4W�z����P   P   Z��9~���ۿ1�F��~���+�CJA�fLR�uPA��5�E�����F�K�ۿN~�v�+3���u�ߗN���t�4'��P   P   �߾R�6�������0�i��#���+�M�0�.�0�S@��S��G<j�������67�I�߾@V���Y�
�Y�];��P   P   F?��{���N��X�0�i��~��XH����Bm��h����Vj�����1���?O��8�dw��u�XY���t�P   P   פ��7`���K��W����0�F��������������#G�����A��l]X�}��,���Ҋ�,�l�c�l�P   P   #Y��N���o�¾�K���N������ۿ���8�6�%E�'7�f���ܿ�D���cO�����þ�畾Vt����z�P   P    B������N���7`��{�Q�6��9~��%��M	Ͽ"�翎��[@Ͽ#j����~�=^7�x[��л��Oч�L��P   P   !����YLپ���?��e/Ծ[����-�\�T��q��g|�F�q���T�7G.�! ���ԾUa���!���Iپ��P   P   ��z��T߾մ�\����������+�Ӿ7��j���"���"�������Ծs ���e������_Ѵ��=߾P   P   �Iپ��B]پ*ᴾ�4��P�p�"�l�z����ޟ��(����Ͼ�-׾X�Ͼ�u��t@��`^��,dm��Xq��?��_Ѵ�P   P   �!���YѾ�^Ѿ�'�������q�unL�*HE��U�PIp��z��g���b���Ⰵ���p�<�U�^�E��L��Xq�����P   P   Va��fFҾ")ݾG<Ҿ�E���/����l��=E�wG3�K�1�|�8�|A�7�D�jUA��z9��2��4�_�E�.dm��e��P   P   ��ԾT���O��G�m����UԾ�����녾��T��1�˜��6������n��(C��2�>�U�b^��u ��P   P   # ���%���;��D���;�L%�g���xӾ����V�o�c�8������f������o���z9���p�w@��ԾP   P   :G.��	_�����Q򒿨䒿6e����^���-��o��Һ��,���@�O7�R���f������mUA�䰅��u�����P   P   ��T�`��������ܿ�x鿧�ۿ����Mi���DT��&�kϾ�-����C�O7������:�D�e���[�Ͼ���P   P   J�q�>M������7	�8���7�G��s{���񮿔q��;"�u�־�-���@����6�A�h����-׾��"�P   P   �g|�!6¿+:�n�T��}��ʩ���a��LET�~��������{��;"�jϾ�,��b�8�̜�}�8��z����Ͼ��"�P   P   �q��&¿� �ʬy�E���g��V��q����Qy���������q��&��Һ�U�o��1�L�1�RIp��(��j�P   P   ^�T��$���!���y�5>�������������Qy�~�����DT��o�������T�xG3��U��ޟ�9��P   P   ��-�m|������`T�-ѳ�����������p���KET�q{��Li����-��xӾ�녾�=E�*HE�z���,�ӾP   P   \��w�^���������Z���M�����������V���a��E��������^�f��������l�unL�#�l�����P   P   f/Ծ�,%�uK��Юۿ��7������M�������g��ȩ����7���ۿ5e��L%��UԾ�/���q�P�p����P   P   @�������c;�_���D+鿄�7��Z��,ѳ�3>��B���}�� 8��x鿦䒿��;�j����E�������4��\���P   P   �����Ѿ]��C�_���Ϯۿ����`T���y�Ǭy�j�T�5	��ܿO��D��G�E<Ҿ�'��)ᴾմ�P   P   YLپ�4Ѿn�ܾ\��c;�uK������}����!�� �):���������������;��O� )ݾ�^ѾA]پT߾P   P   ������4Ѿ��Ѿ�����,%�v�^�l|���$���&¿6¿;M��]����	_���%�Q��dFҾ�YѾ��z��P   P   ���x���kG�/3�9pھ� ϾDJ��`0�iG�9~O��G�֐0�������aiϾ��ھ"�)�F�V{��P   P   V{��t����SV�wP��վ;{��de���뷾�۾K{��U��F��
���q,ܾ�D������㕥�G�վ�#�V�P   P   )�F�e?Z� G��U�\4׾k��8Lr��fr�|)��W*������j2��z����i��Xv����r�ԣr�	����־�#�P   P   "��t&�ʃ&��C��վN$��?�Z���9�6�;��P�P*h��w��>w���h��Q�se<��:�\[�	��H�վP   P   ��ھb����������ھ�����Pr�7�9������w�#�yi,�070���,�D$�H���d ��:�֣r�䕥�P   P   ciϾF[��G��D�)I��,AϾ�g��pEr�<�;����j����F��g�4	����I��ue<���r�����P   P   ������C'�/��.'��l�XJ�]̷�����`/P��C#�C��L������/��4	�F$��Q�Zv���D��P   P   ���.�:���^���s���s�O^�ʘ:�6��3�۾$ٟ�d�g���+���������g���,��h��i��u,ܾP   P   ِ0�Pl�eؔ�X���׶��8�������k��&0� ��	'��|Zv�O�/����M���F�270��>w�|������P   P   �G�ы��ᱽ����N� B�L_�1e��E��D�F��p�]���|Zv���+�D�����{i,��w�m2��H��P   P   <~O��(��?�޿���=�8M�(o=��P��o޿ޙ��O��p�	'��c�g��C#��j�y�#�R*h�����W��P   P   kG�>��r�뿻�.��4o�����6����n��J.�XT�ޙ�C�F� ��#ٟ�_/P������P�X*��N{��P   P   `0��o����޿My.����X���$���E���ǁ��J.��o޿E���&0�2�۾����;�;����7�;�})���۾P   P   ��� �k������f�|o�DS��c���]���E���n��P�/e���k�5��\̷�oEr�7�9���9��fr��뷾P   P   EJ��:�����_��m=�₎��#��c���$��4���&o=�J_���ɘ:�VJ��g���Pr�?�Z�9Lr�ee��P   P   � Ͼ�V�)/^�I ���.���L�₎�CS���X������5M�B��8��
O^��l�*AϾ����N$��k��;{��P   P   9pھ�	��6'���s�֨���.��m=�zo� ���4o��=��N��׶���s��.'�'I����ھ�վ\4׾�վP   P   /3��������.���s�H ��_f�Ky.���.�|����X����s�/��D����C��U�wP�P   P   kG�y&�w����5'�(/^����������޿o��;�޿ޱ��cؔ���^��C'�G����Ƀ&� G��SV�P   P   x����NZ�y&�����	���V��:���k��o��<���(��΋��Ll�+�:���C[��a���t&�e?Z�t���P   P   +�����<=���ih��V�J�־�eѾqg��#�f��H$�a��"F�C��ƦѾ��־<A�&h����Y��P   P   Y������jϿ����X|"�A˾����m��h$����Ͼ�߾�߾/�Ͼb��Z���!"��˾�9"�]��o*ϿP   P   �����п�<��������+�Ib;p1��Ghc��(o�����6"��Û�M>���燾��o���c�1+��l;O0+�]��P   P   &h��f���z��jh��"��m;'&��s;�8c+��t8�>M���Z�[�[M���8���+��L;����m;�9"�P   P   =A��k6��(F� �6�`q��]˾�6���
;����*�����l"�r�&��T"�<9����q��L;�2+��˾P   P   ��־������*�������־U��Kc��9+�_z�C��\'�o|	�]�	�b|��(�����+���c�#"��P   P   ɦѾ+����<��t��ط��dѾ�P����n�#8�e��K�<* �����i �b|�=9���8���o�\���P   P   G��+��l4��XE��KE�H4�����7�ߵ�9l���L��!��4	�>������^�	��T"�[M��燾b��P   P   $F�59�	'e�Q���r���=x����d��8����u-Ͼ����BGZ���%��4	�=* �p|	�s�&�[�O>��3�ϾP   P   d��wX��S��TL���ſ�ᵿ�X#��,���X�C����޾sG��BGZ��!�K�\'�m"���Z�Û��߾P   P   H$�dgk��\��V�ӿ����?�������mӿ�����j���#���޾�����L�d��C�����@M�7"���߾P   P   h���Yk��c����V[��W/��K/��=�@쿱&����j�C��u-Ͼ9l��"8�_z�*���t8�����ϾP   P   �#��RX��K��~y�J�"�u�J���[���J�A�"�@쿸���X����ߵ���n��9+����9c+��(o�i$��P   P   sg�m�8�o7��j�ӿP�W�J�
�m�<�m���J��=��mӿ+���8��7�P��Kc��
;�t;�Hhc��m��P   P   �eѾv��I�d��(�����N/���[�	�m���[��K/�����V#����d�����dѾT���6��'&��p1�����P   P   K�־���@44��k���������N/�V�J�t�J��W/�>��ߵ��<x��H4�׷���־�]˾�m;Jb;A˾P   P   �V�Z��J��
!E�`㉿�������P�I�"�T[������ſ�p����KE�s�����_q��"���+�X|"�P   P   �ih�t6�������
!E��k���(��h�ӿ|y���T�ӿQL��O����XE�;��)�� �6�jh���������P   P   <=��&y��cF����J��@44�H�d�n7���K���c���\���S��'e��l4�������(F��z���<���jϿP   P   ��� ѿ&y��t6�Z�����u��l�8��RX��Yk�agk�wX�29��+�*������k6��f����п���P   P   E}��Oj��K$�=.��³F�������þ+�ݾW���"������}�ݾE�þx ���x�UxF��뻿_$�7.j�P   P   7.j��Fj�?�8�{r�7�w�cq��襾�,�����é��%���1���㩾՗�mI���٥��;�(Ww�� �j8�P   P   _$�4#9��L$��z�����Tݡ�Lyd�kX�(�m�L�����Lׂ���m�[�X���d�j���������� �P   P   �뻿����EB��;�w���֜��W7N��y*�}0��BC���P��Q��}C�f�0�д*��&N�[H����)Ww�P   P   UxF�l?���퐿�f����F� ���顾2N��F�����غ+��41�Y�+���9p����&N�k����;�P   P   �x�k���5�y�5�O�����0���)dd�lT*�#��h����s� ��� �v���}�:p�Ҵ*���d��٥�P   P   z ���񾓗�#�����
��������X��+0�9~��h��������w����h�0�^�X�oI��P   P   H�þ8p��o4�������6��*���aþ�n���$m�*�B��V+�͒ �&������ �Z�+��}C���m�!՗�P   P   ��ݾ���|�+��C�ĭK�g�B���+�gG��dݾMc��(e��vKP�K�0�͒ ����t� ��41��Q�Nׂ��㩾P   P   ����B"�9OM� �s�{�������=�s�M���!��(��$����5��vKP��V+��h����غ+���P������1��P   P   %���A+/���g�|����ק�3���k���9א���g���.��j��$���(e��*�B�8~�h�����BC�M��%��P   P   Y����"/�8�q�*���-ÿ>ڿ��ٿ�ÿ�垿�q���.��(��Lc���$m��+0�"���}0�*�m��é�P   P   -�ݾ,,"���g��	��:�Ϳ/����-��ܚͿ�垿��g���!��dݾ�n���X�kT*��F��y*�kX�ﬗ�P   P   ��þ�e�5.M��퐿�#ÿh,���	�z�	�-���ÿ8א�M�gG��aþ���(dd�2N�W7N�Myd��,��P   P   ����3����+�a�s��ȧ���ٿҰ��	�����ٿj���<�s���+��*�����/����顾ל��Uݡ��襾P   P   ������B�	���������ٿg,��/��=ڿ2�������e�B�5����� ������cq�P   P   ³F��k�vz������K�����ȧ��#ÿ9�Ϳ�-ÿ�ק�y���­K�������N����F�;�w���8�w�P   P   =.���P����5�3�����
�B�`�s��퐿�	��(��z�����s��C����"��x�5��f��FB���z�|r�P   P   �K$���琿��5�vz�����+�3.M���g�6�q���g�7OM�z�+�m4������5��퐿뿮L$�?�8�P   P   Oj�469��뿁P���k����3���e�*,"��"/�?+/��B"����4p����k�l?�����5#9��Fj�P   P   �7�������y�j�
�������ޱ����V��������ǾS���l-������s߱�����焿�~
��y����P   P   ������Ћ�%�.��°���'��'��lE��5��������h��[+��n���1I������h'��Z��J_.�ީ��P   P   �y�����y�$�.�2�ÿ�A�SMž�'w�ՏV��d��?y�-+��	]y��Id�/�V���v�&�ľ��@�9cÿJ_.�P   P   �~
�ɺ/��/��
�qܰ���A�n0;/s��`>��@�!�T�o�c�)�c���T��A��r>�%�r��̾��@��Z��P   P   �焿�o���Fʿ֭���:����'��bžs���7��m1���A�VT�Dg[��(T��7B�S�1���7�&�r�&�ľ�h'�P   P   ���w�7���Y��Z��>8�4��B��1w��=>��S1��O<��M��Y��Z��-N�Y�<�S�1��r>���v����P   P   u߱����M�	�K����	���澴��2��GGV�u�@�ݹA���M��Z��_�(=Z��-N��7B��A�2�V�2I��P   P   �����Ⱦ��뾟%�B#���뾿�Ǿ�Z��FY����c��$T��S�0�Y�s�^��_��Z��(T���T��Id�p���P   P   n-��e׾���X��4�����)���'�־�ů�Ӿ��7�x�m�b���Z�/�Y��Z��Y�Eg[�+�c�]y�]+��P   P   U����/���GF*��&8��8��"*�6��ط�[h����ƀ�m�b��S���M��M�VT�p�c�.+��j��P   P   ��Ǿ�[���#�E�G_���h��*_�<lE�Do#���GǾ�7�x��$T�ݹA��O<���A�!�T��?y����P   P   �����V��*�{FV�z�}�%���׉���_}�6V���)��Zh��Ҿ����c�t�@��S1��m1��@��d���P   P   W�����#�AV��u���旿�G���ڗ�(a��5V�Do#�׷��ů�EY��FGV��=>���7��`>�֏V�6���P   P   �����־-��P�E��}�j旿�.��c*���ڗ��_}�;lE�5��&�־�Z���2��0w�s�/s��'w�lE��P   P   �ޱ��Ǿ�����1*�:_�֏��9K���.���G��։���*_��"*�'�����Ǿ���B���bžn0;SMž�'��P   P   �����;�����8�2�h�֏��j旿�旿$�����h��8������뾢��4���'���A��A���'�P   P   ���m8�$�	��
� ���8�:_��}��u��x�}�G_�&8�3��A#���	��>8��:��rܰ�3�ÿ�°�P   P   j�
������Y����
����1*�N�E�AV�yFV���E�EF*�V���%�J���Z�֭���
�$�.�%�.�P   P   ��y�{�/��8ʿ��Y�$�	�:�뾭���,���#��*���#����������L�	���Y��Fʿ�/���y�Ћ�P   P   ���J���{�/����l8�����Ǿ��־��V��[��/�b׾�Ⱦ���w�7��o��ɺ/������P   P   ������Ѳ���v1�����W������򩎾�����T��xϥ��]�����^����v�����)Q���?1�G�������P   P   ����b�������~�`�O�޿��G���Ⱦ����D�"^��<���@���h���T�8���Ⱦ�dG�w!޿l�`��֭�P   P   F������������`�����B�m���辄̌�(nn��z��r���J��|��$�z�umn����r%��m�7��l�`�P   P   �?1�)Oa�wra��1���޿��m�>���H���8k���q�ҷ��"��0(��ǅ���q��+k�e���
���m�w!޿P   P   )Q�����������𻢿�H���������k���o�?���ԓ�2��䓾)X��!�o��~k�f���r%��dG�P   P   ���_�O�F�y���y�Y	P��
�[!ɾSɌ��k���o�vΆ��g��`ȡ��ҡ�5�������"�o��+k�����ȾP   P   �v��4�ྪ~��������O���� ���#n�saq�����V�����>P���.��5���)X����q�vmn�9��P   P   _����姾=5þS;վ/=վ�4þԧ�,�����~��,z��x������|����A��>P���ҡ�䓾ǅ�&�z��T�P   P   ���Y?�������о(ؾ�о3㽾W���m���(�����+Ԏ�$���|������`ȡ�2��1(��|���h��P   P   �]��v,����Ҿ�K쾟���ڟ��j�x}Ҿ�ȶ���ӑ��茾+Ԏ������V���g���ԓ�"���J���@��P   P   yϥ��xþQ��k��D��l��0��F�x��|
þ`���ӑ�����x�����uΆ�?��ѷ���r��<��P   P   �T���sþW�𾼰���%��x2��n2���%����?.�|
þ�(���,z�qaq���o���o���q��z�"^��P   P   �������h辈��K�,��PA���H��?A��z,����w���ȶ�l�����~��#n��k��k��8k�(nn��D�P   P   򩎾�-��ѺҾ�e���%��QA�cQ��\Q��?A���%��F�w}ҾV���+���� ��SɌ����H���̌����P   P   �����ק������9�-A��{2��I�cQ���H��n2��0�i�2㽾ԧ�O���[!ɾ���>���¶���ȾP   P   W��\���þ��о�����p��{2��QA��PA��x2��l�؟���о�4þ��ྸ
��H���m�C�m���G�P   P   ����ҼO�Pk��վe�׾����,A���%�J�,���%��D�����&ؾ.=վ���Y	P�񻢿��޿����P�޿P   P   �v1����<y�����վ��о�9��e��������k��K쾻�оR;վ���y����1���`�~�`�P   P   Ѳ��aa�����<y�Pk��þ����кҾg�U��O辩�Ҿ���;5þ�~�G�y�����xra���������P   P   ���!��aa����ҼO�[�ྯק��-������sþ�xþt,��W?���姾3��_�O����*Oa����b���P   P   ����z����̫@��'�����"����$�������v���s��y��ݠ��E���z��מ��󭿬z@����jn��P   P   jn��Oy��!:���<t�����W�L�׾?��UǊ� r��������t��-Ċ�g%��O�׾��V�@��s�?��P   P   ����.�����Lt�zo�z���C�Z���6&���|��1ܪ��谾rા���%���r���� �������s�P   P   �z@��t��6t���@����)���gF
�����ᥚ��Ͽ���%Ǿ�)Ǿvɹ�%�������PJ��6�	����@�P   P   �󭿷G��V�����c���HW�S�?����J���l����žX�۾A��2�۾FƾA|��?��PJ���� ���V�P   P   מ��V��V���l���/W����n"ؾZ���я��\��^�ʾ���F���P��p�羝�ʾA|�������r��P�׾P   P   �z��԰׾`��
��,��׾����>)������A���p�ž���[� ��T�ť �p��Fƾ%���&��g%��P   P   F�����CM���*���/���S������h�������j1��aw��E[۾� ��)L��T��P��1�۾vɹ����-Ċ�P   P   ޠ��}���đ�(��mŝ��������~T��AO����{����ƾJ��� ��[� ��F��@�㾡)Ǿrા�t��P   P   y��&7�����X��y«�ͳ���,��=Ǜ��ڔ����r����~����ƾD[۾�����W�۾�%Ǿ�谾���P   P   �s������^������/ž��ɾ�ž'Ѹ�W���W��|��r���{��`w��o�ž]�ʾ��žϿ��1ܪ���P   P   �v�������c��Lfƾp�ھ����澊yھ�ƾ���W�������i1��@���\���l����|��r��P   P   ����m3���\��fƾh��H)��� �[��ߦ⾨ƾW���ڔ�@O����������Џ���J��ग़�5&��TǊ�P   P   �$�����I��E���ھ�-�����ޱ�[���yھ'Ѹ�<Ǜ�}T��g���=)��Z���?�������Z���?��P   P   "����������T���5ž���� ����� ��澿ž�,��������������o"ؾS�hF
��C�L�׾P   P   ���,�׾�;������ū���ɾ����-��G)����澫�ɾ̳������S���׾����HW�)���z���W�P   P   �'��R�V�Z� �c��Ƽ���ū��5ž�ھg��o�ھ�/žx«�lŝ��/���,��/W��c�����{o����P   P   ͫ@�3R��>��]�	�c������T��D��fƾKfƾ���X��(���*���
��l�������@�Lt��<t�P   P   ��\t�@��>��Z� ��;������H���\���c���^�����đ�BM��`��V���V��6t����":��P   P   �z���1��\t�3R�R�V�+�׾�����l3���������%7��|�����Ӱ׾�V��G�t��.��Oy��P   P   �v��f���k5��c�0�g��G���{���ю�
;��i������0����3�����[��n�1᡿_�0��#���y��P   P   �y��q��������`�_J࿹oO����E)������k���J�þ0�þ����=�������R�*O���߿�e`�H|��P   P   �#���v���?��D�`�PD��^@y�H���þ�����~Ӿm�辸l�����yӾ)����Vþ�;�	�x�s����e`�P   P   ^�0���_��`�0�0�fv࿯Xy���F�վ9pѾU*�4���E��F�z��D*�0\ѾSվM���x���߿P   P   0᡿��ݿ����#�ݿ�A��v�O�|��g�վ&�ؾC��������&��[-�*�&�e������o�ؾSվ�;�*O�P   P   n��G���l���l�&qG����ڼ��|þ�PѾ����)��?3�Q0B��5B�O3��"�����0\Ѿ�Vþ�R�P   P   �[��jyȾc�羀��h'� �Ⱦ����p�� a�����r��23�A�I��[R���I�O3�e��D*�)������P   P   ���懾�n��*���􍒾�q���؇�����N���Ӿ.��؂&��B��PR��[R��5B�*�&�z���yӾ=���P   P   �3���-���m�n}j�i�j��Zj�N�m�`�~��ړ�1���k辵��--��B�A�I�Q0B��[-��F���辟���P   P   0���E[��+Az�m�p���n���n���p���y�������{þ���؂&�23��?3���&��E��l�0�þP   P   ���"9���7���P��P���qB���������y݇�xȑ�֏���{þ�k�.��q��(����3��k��I�þP   P   h����:�����Ȳ��BB���Ö�B���	��0g��਌�xȑ���1���Ӿ������A���S*�~Ӿj���P   P   	;��`���;��嵎��������Y�������_��0g��y݇�����ړ��N��a���PѾ%�ؾ8pѾ��������P   P   �ю�a<�cNz�;Y���K����8���.}������	�������y�_�~����p���|þf�վE�վ
�þD)��P   P   �{��\��m�4q��̅�aז�m��8����Y��A���������p�M�m��؇�����ۼ�|����H�����P   P   G���Ⱦ�g���j�co��_��aז�
�����Ö�qB����n��Zj��q�� �Ⱦ���x�O��Xy�`@y��oO�P   P   h���G�M��Ns����j�co��̅��K������AB��O�����n�h�j�󍒾i'�'qG��A��hv�QD��`J�P   P   d�0��ݿ
�l�����Ns���j�4q�;Y��嵎�Ȳ���P��k�p�m}j�*��������l�%�ݿ2�0�E�`��`�P   P   l5����_����
�l�M���g����m�cNz��;������7��*Az���m��n��c�羦�l������`��?������P   P   f���v����_��ݿ�G��Ⱦ\b<�`���:��"9��E[���-��懾iyȾ�G���ݿ��_��v��r���P   P   EL���)���x���	��S��Q���ڱ��բ��)V���=Ⱦ�L��Fz������=���q��t<��1�	���w�`#��P   P   _#��#+��p����.�򈴿.p7�����gȾg�׾�����g�����P�׾fAȾxF�|,7�F���r.�����P   P   ��w�ߊ�Ix�ʴ.�0ɿMAY���	�9V쾥����w�D$��*��@$�p����!���	���X���ȿ�r.�P   P   0�	��b-�]y-��	�b���jRY�Q��?X��=���*�acF�K&W�&W��bF�7�*�x2�Z:�t����X�F��P   P   s<��A����¿-���Հ���7�:�	��Q���8�O.`�ɞ~�����~��6`��8����Z:���	�|,7�P   P   q����&�\@�v@�'���r�澖0�j%��8���i�i,��Κ��{���'6����i��8�x2�!�xF�P   P   =���5���(eľ�-̾��ľC���ZƱ��(Ⱦ=o����*��`�^!��B��<������'6���6`�7�*����fAȾP   P   ����d/���v��#r��#r�Yqv����a���>׾�4�MF��c~�f���5���;���z�����~��bF�p�P�׾P   P   Fz��Q����YV�p�=�t�6�&�=���U�Gc��n��R���#�U�V��ꄿf���B��Κ����&W��@$����P   P   �L���F���d�@���0���0�_$@�2oc��א�=����o�Fa*�U�V��c~�]!��h,��Ȟ~�J&W��*�g��P   P   �=Ⱦ�7���6y��@T�~eA���;�� A�ԷS�mx�����Ǿ�o���#�LF��`���i�M.`�_cF�D$����P   P   (V��b<���$���.c�aS�0+M��M���R� �b�M������=���R��4���*��8�	�8���*��w����P   P   싰�%T��EJy��:c�%�Z��Y�$Y���X�n>Z� �b�mx��א�m��>׾;o��i%� ��=�����e�׾P   P   �բ�.��.d��aT�X~S��.Y��^��^���X���R�ӷS�1oc�Gc��`����(Ⱦ�0��Q�>X�8V��gȾP   P   �ڱ�+C��Y}V���@�C�A�WaM��RY��^�$Y��M�� A�_$@���U����YƱ�q��:�	�Q����	����P   P   Q��������v�C>�n#1��;�WaM��.Y��Y�0+M���;���0�%�=�Yqv�C������7�kRY�NAY�.p7�P   P   �S��@�&��Lľ�r�!7�n#1�C�A�X~S�%�Z�aS�}eA���0�s�6��#r���ľ'�ր��d���0ɿ󈴿P   P   ��	��z��/@���˾�r�D>���@��aT��:c��.c��@T�@�o�=��#r��-̾�v@�.����	�˴.���.�P   P   �x�bX-��b¿/@��Lľ��v�Z}V��.d�FJy��$���6y��d��YV��v�(eľ\@��¿^y-�Jx�p��P   P   �)��(ڊ�bX-��z��@�&�����,C��.�&T��c<���7���F��Q���d/��5�����&�B����b-�ߊ�#+��P   P   �0����g��"��^���KE�8�쾊&��Dľfr޾	e��b����T��aT޾��þ����2���/E�&M��i�"�G�g�P   P   G�g���g��J7�K���W�����R���������_�"�޺/�t�/���"�U��������G���0�����}/7�P   P   i�"��6��"�G�迋ۏ���4�}��t�l,���M�?�h���r�>�h���M�&X,�FY��Q���4��������P   P   &M����{&���l����4�X������C�-�t�G���嵟�����/�����t��C����lz���4��0��P   P   �/E��u�U܅���u��~E����v� ��@L����ބ���
Ŀ`�ο;Ŀ����E��`AL�����Q�G��P   P   2��S�����B �%�������S��mC�+���]��oۿ\c��i��)ۿAp��E���C�EY����P   P   ����ki���������0���t���켾S��x*,��rt�5d��_�ڿES��
�>^�)ۿ������t�&X,����P   P   ��þM5��d��wM�amM���c������þ̖���M��U��i�ÿ4=��H�
��
�i��:Ŀ/�����M�U��P   P   `T޾+𗾫wX�9*�.���*�[X�Б����ݾ%Z"��4h�au��@uο4=��ES�[c��_�ο����<�h���"�P   P   �T��3����m��j0���-��A 0��4m� ���T����H/�*Ir�au��i�ÿ^�ڿnۿ�
Ŀ䵟���r�s�/�P   P   `�������肾T;C�g�����4���B�,s��굾����H/��4h��U��4d���]��݄��F���=�h�ݺ/�P   P   e��⏶��ɇ���P��w+�X(����+��%P�E��굾T���$Z"���M��rt�*�����+�t���M�^�"�P   P   dr޾�5��z��� �P���0��f �VO�> ��\0��%P�,s��������ݾ˖�w*,��mC��@L��C�l,����P   P   Bľ��=$n�AlC�e�+��~ ��|�_\�> ��+���B��4m�Б����þQ���S� ����t�����P   P   �&��.W��θX���0�Q��am�0���|�VO����4�A 0�ZX�����켾��v�W��}�Q��P   P   7��e����5d��~*��1��)�am��~ ��f �X(���,���*���c��t���������4���4����P   P   �KE������ޛM�>��1�Q��e�+���0��w+�g����.��amM�0��&���~E��l���ۏ��W��P   P   �^���u�C��R���ޛM��~*���0�ClC�"�P���P�U;C��j0�9*��wM�����B ���u�����I��L��P   P   �"����8���C������5d�иX�?$n�{����ɇ��肾��m��wX�d�������V܅�}&��"��J7�P   P   ��g�;�6�����u���e���/W��	���5��䏶����4��+�M5��li��T��	�u����6���g�P   P   ���+ �ָ�,�e��X� h־��Ѿ�+�K���g��$��Z�l�����x�Ѿ�1־�A�>�e��ϸ��) �P   P   �) �$/ �Tο^苿F5��4�����t�g�9�rY�@l��l�w Y�r9��S�+��-���4�=͋�S;οP   P   �ϸ�г̿�鸿��f�D�8%�(���4�7�e�!č�nꢿ� ��i⢿����3�e�՝4�M��R���`D�=͋�P   P   =�e���Q����f��)5��$�ʨ�I�E��烿ެ�ywԿ>~�z�nԿӬ�M܃�R�E�L��R����4�P   P   �A��� ���)��!�0j�b0�c����E�O[���j������
�*�#�w�) ���l���[��R�E�M��-�P   P   1־� ʾ�˾��˾# ʾXJ־|��o�4�\˃��T��.D� -0�L�K�<�K�890�R��l��M܃�՝4�+��P   P   w�ѾȺ��ʗ���n��▆�魝�4aѾ�+�ce�����v���d0��\�pLo���\�890�) ��Ӭ�3�e��S�P   P   ���"����8c�C�:��:���b��W���� 9��{��Կ�����K��9o�pLo�<�K�w��nԿ����r9�P   P   k��X���po�]+�����+���n����'/�@�X�Ύ����AM#���K��\�K�K�)�#��z�h⢿u Y�P   P   �Z�Yо��Ŝ8����3j�� 8�����vϾO���k�񟪿�����c0�-0�	�<~� ���l�P   P   �$���\g��qEM�c�������ȒL��ܕ��B߾Q:$��k�Ύ��Կt���-D�����wwԿlꢿ>l�P   P   �g�R����O0[��"��O��h�!�SZ�<k���B߾O��?�X��{�������T���j��ެ� č�pY�P   P   J��18оI}��VG[��&� U	������	���%�SZ��ܕ�vϾ'/� 9�ce�\˃�N[���烿4�e�e�9�P   P   �+񾕶��'��e�M�RO"��q	�~���E���	�h�!�ȒL�����������+�n�4���E�G�E��4��t�P   P   ��Ѿ�˟�l�o�v�8��5��[�F5 ��������P����� 8���n��W��3aѾ|��b��ɨ�'�����P   P   �g־�松��c��+������[��q	� U	�����3j��+���b�魝�WJ־b0��$�7%��4�P   P   �X�ʾ*���I�:��X����5�TO"��&��"�d���������:�▆�# ʾ0j��)5�g�D�F5�P   P   -�e�s� ���˾"���J�:���+�w�8�g�M�XG[�P0[�rEM�Ɯ8�	]+�B�:��n����˾�!��f���_苿P   P   ָ��冿n�)���˾*�����c�o�o�)��J}�����]g����po��8c�ʗ�� �˾��)�R����鸿TοP   P   �+ ���̿�冿s� �ʾ�松�˟�����38оT���ZоY���#���Ⱥ��� ʾ�� ���ѳ̿$/ �P   P   ؊���=�,~D�����\پ2 Ͼ5��N'�*�0�?�G���O�EG�3�0�����V�ξ&پ����tD��:�P   P   �:��C�_W��$�&��T���7���6;���l��挿;��������Ռ��gl��;��}�4���@��h�$�HW�P   P   �tD�'VS��D�z�$����f�
�tR'�D�^��1��:��X�߿�z�s߿�!��G����^��''��
�+��g�$�P   P   ���t������7��U�
�9/�4Zt������V��_7/�3/���a?�̬���6t�5�.��
�@��P   P   &پ�Ӿ
վ��Ӿ9Mپ���/4'�?t�qD�����L>��Gp�e���6Ep��I>�����@���6t��''�4���P   P   V�ξr����������Ĥ���ξ@s���^�͗�����M��6��v2��86��1@��6�M����ˬ����^��}�P   P   ���P����q�P�Y��q�[3���\�\�:�f픿,�>��#�����Xp��� ��1@���I>�`?�F���;�P   P   ���2��zr�jZ9�1@9�&r��ⷾ����k��ν�A����o����q_��Wp��76��4Ep����!���gl�P   P   2�0�9Nܾ�b��7�;����H�;�8��O�۾e0�΄����޿��.�{M��������u2��d���3/�	s߿�Ռ�P   P   DG�C
���x���P��>����NP����K��!�F��&���뿨�.���o��#���6���Gp�]7/��z�􍚿P   P   ��O��	��ﱾ�h��#�G|��S#�r�g��O��ʙ�J\O��&����޿@���>��M��L>��V�߿:���P   P   =�G�p	�����Eyw�j�,�f�����>�+��}v�vѷ�ʙ�!�F�̈́���ν�*�������V� :���挿P   P   (�0��6��3����w�#\0�GK�7���M��̣/��}v��O��K��e0��k�e픿̗��oD�������1����l�P   P   L'���ܾ�����h�C�,��l����Dm�M��>�+�q�g����N�۾���[�:���^�
?t�2Zt�B�^��6;�P   P   2��Gz��ѣ��TQ�%$�O?	�$�����8�������S#��NP�7���ⷾ�\�?s�.4'�8/�rR'�6��P   P   0 Ͼ��� s��<������P?	��l�HK�g��H|���G�;�&r�Z3����ξ���U�
�e�
�R���P   P   �\پ�,r�l�9��s ���� %$�D�,�%\0�k�,���#��>����0@9��q��Ĥ�9Mپ7�����%��P   P   ���&�Ӿ*4��fLZ�m�9��<�TQ���h���w�Hyw��h� �P�7�;�jZ9�P�Y������Ӿ���z�$��$�P   P   -~D��q��վ*4��-r� s�ң�����4������ ��x���b��	zr���q����
վ���D�_W�P   P   �=��KS��q�'�Ӿ����Iz����ܾ�6��r	��	�E
��:Nܾ�2���P��r����Ӿ�t�'VS��C�P   P   �.���_�־Э��������Ծ����.�� U��r�m�|��r���T� R.����.ԾLw��|��&�־*{��P   P   *{��3���q��3�Ͼ<_Ѿ/����%�hZ_�n�,���	�¿U�¿�����ѐ��_��g%�X|��@Ѿ�SϾA��P   P   &�־Ofܾ��־�Ͼ� ܾ4$���;�^����O���v����� ��+���M��(&�������;����۾�SϾP   P   |��精-�4����FѾ��"D��"��\qܿ�n��;U�`�z�T�z�1&U��W��Kܿ���J�C���@ѾP   P   Lw��5��7��m��� �������;�������̈8����Ȓ����������}8���������;�W|��P   P   .ԾGÓ�E�o�a�o�f���k"Ծ�Y%������6ܿm8�"���-���9��;�@8���-���}8��Kܿ����g%�P   P   ���#ͪ��l�'L�j`l�l���w��G�^�����+��ĉ�����y� w����?8�����W�'&���_�P   P   �Q.���Ӿ���IOE��0E��셾*�Ӿ�.�����������T�YI��T�Vk� w��;����/&U��M���ѐ�P   P   ��T����p!���KU��h3���T��Ɵ����ywT�f)��09���y�����S��y��9���R�z�*������P   P   �r����"{��Y�p��2���1��p�$�kD�_Wq�e¿�)���y�YI������-��ƒ��]�z����T�¿P   P   j�|��"���Ͼ���I09�ɿ���8��?��9Ͼ�["��!|�e¿/9���T��ĉ�"������;U�����¿P   P   �r�j�"�L�׾�ɍ�3HA�_U�� �B�@�@?����־�["�_Wq�e)�������+� m8�ʈ8��n��v��*���P   P   � U���оDڍ�g�D�Ƥ�����@���C�??��9ϾkD�xwT���������6ܿ���Zqܿ�O��l�P   P   ��.���������݅�"�A�%���������@�B�@��?��#�����.�F�^���������"��]���eZ_�P   P   ���HԾ�r��:7q�(�9������������� ���8��p��Ɵ�)�Ӿv���Y%��;��"D���;��%�P   P   ��Ծl$���s���U���2�m����&��Ǥ�_U�ɿ���1���T��셾k���j"Ծ����3$�-���P   P   ��������$m�5F��64���2�)�9�$�A�i�D�5HA�K09��2��h3��0E�i`l�e��������FѾ� ܾ:_ѾP   P   Э��󲖾j^p��L�6F�!�U�<7q��݅�Fڍ��ɍ����Z�p��KU�IOE�'L�`�o�m���4����Ͼ2�ϾP   P   _�־Y���.��j^p��$m��s���r������оN�׾��Ͼ${��q!������l�E�o�7��-󲾚�־q��P   P   .���oܾY���������n$���HԾ���!��l�"��"���������Ӿ#ͪ�HÓ�5��精Ofܾ3���P   P   � ��㪃��I��Q7���b��n�ʉ��[F�V�t�ċ��O��~���Jgt��F�UG���߾�������!��ŗ��P   P   ŗ������}w������_��~P��w7���~�K���M�Ͽj迤��jϿ�q��ƣ~�/7������Ӕ��U��P   P   !��7x�l7��������¾��2yO��f��(Jܿ�1��{7��E�qf7���Eܿ�7���4O�3W�W¾Ӕ�P   P   �����j���j�����9���y�#mX�(c�����VZG�hd��td���\���Q���2G����;��:X�3W����P   P   ����s�e�W�)t�B���$�<JO��M�����j����� ��rn�r���	����j�����;���4O���P   P   ��߾:&���Y�Y�!��5�߾�$7�
/������j�P������1�)1����������j����7��/7�P   P   TG�{Q���u��yN�Q�t��*��/%�/i~�e�ۿ��F�w޶�}�j�A���R��A����	���2G�Dܿţ~�P   P   �F��g�[8���WW��8W�G������E��,�����r�����A�0��R���R�)1�q����Q�����q��P   P   Hgt��|n��$�o�p�I���o������4�s�6�ο��6������8�@�0�i�A��1�qn��\��of7��jϿP   P   }����J+���Ӿ�臾�~I�;LI�����#AӾ��*�S���]�"�D��������}���� ��rd���E���P   P   �O���b9����v��{xP��2��	P�������S�8��ݑ��]翘�6�r��u޶�N������fd���{7�g�P   P   }ċ��o9��*�A��LX��'��'��uW�h����L�S�8� S��5�ο�����F��j��j�SZG��1�J�ϿP   P   T�t��m+��꾧/���a[��#�:w�0#���Z�h��������*�3�s��,��c�ۿ��������&JܿI���P   P   �[F�JB��Ծ����[fX���#��
�r
�0#��uW����"AӾ����E�-i~�	/��~M��&c���f����~�P   P   ɉ�J��{δ�:���Q�!0(�����
�:w��'��	P����������.%��$7�:JO�!mX�0yO��w7�P   P   k�ܽ��!���h�p�=AJ���3�"0(���#���#��'��2�:LI���o�F���*��3�߾�$��y���|P�P   P   �b��g�����u��-X�r�J�>AJ��Q�]fX��a[�NX�|xP��~I�p�I��8W�P�t�!��@���9����¾�_��P   P   P7���t���Y��CO��-X�i�p�:�������/��B��v���臾%�o��WW��yN�Y�(t�����������P   P   �I���>k�wX���Y���u�#���}δ��Ծ���*󾵹꾩�Ӿ}n��[8���u��Y�e�W���j�l7��}w��P   P   㪃��lx��>k��t�h���޽��M��KB��m+��o9��b9��J+���g�|Q��:&���s��j�7x�����P   P   �������"8� "n����6h�!""�V�7���t:���%&��֒����U���!����$*����m�ӻ7����P   P   ���b��5�9�0�x�T^��b���C�U����<��忘� ��� �j�����ٌ��T2C�v������E"x��z9�P   P   ӻ7�0$�y�7�ӄx�j鹾ڏ���\�-��N��o'��Q�hb���P��E'��h�֥�C\�IU�
���E"x�P   P   ��m�+6�W/6��m�1���~���e�����
e�6]c��������,���6����$c�D<��y��ëe�IU�����P   P   $*��/�^�#=���^��@��ͣ��c\�h���H����gi��~�����k��
P���؆� h��y��C\�v��P   P   �������T���T��������/C�7ե��;��؆��E��J,�_VM�eVM�!J,��E���؆�C<��֥�T2C�P   P   ��!��nþxf����V�'W��Mþx�!�}s��m9�R�b�[(�� 6,��:_��Nq�F_�!J,�	P���$c��h�،��P   P   ��U��D��Sg��,�g���g�!9������^|U�o���� '�ó���s��4M��Bq��Nq�dVM�j��4����E'����P   P   Ԓ����hþo}���I\�{S��O�¾*g�/N��oe��yP������R��4M��:_�^VM����*�����P�h��P   P   #&��C9��侇���:�\�9]\�d���S侟�8������v �6�a������s��5,�J,�}������hb��� �P   P   ��xH��S��������c��D�\c�t�������b�G�����v ��yP�³��Y(���E��di������Q��� �P   P   r:��2�H�)�� ���k�"�7��w7�=fj�:l��x��b�G�����ne�� '�P�b��؆���3]c�o'��P   P   5����A9�_������Nn�$�2�³�1�2��vm�:l��������8�/N��m���k9��;�F��e�K���<��P   P   V�����4�]5���[k��3�VU��$�1�2�=fj�t����S�*g�\|U�|s��6ե�f�������+��T���P   P   ""�����ـþ�	���d��&8� �VU�³��w7�\c�d��N�¾����v�!��/C��c\���e�~�\��C�P   P   3h�S�þ=۟��肾Z\]�6�D��&8��3�&�2�#�7��D�9]\�{S�� 9��Mþ���̣��~�ُ�`��P   P   �������؀��h��A]�[\]��d��[k��Nn��k���c�;�\��I\���g�&W������@��1��h鹾S^��P   P   �!n��`_��U�,�W� �h��肾�	��_5������ ����������p}��,�g���V���T���^�}�m�фx�.�x�P   P   �"8���6�	�=�	�U��؀�?۟�܀þ�4�a��)��S��	��jþSg��xf���T�"=�V/6�x�7�4�9�P   P   ����Q$���6��`_�����U�þ��������A9�4�H��xH�E9����D���nþ���/�^�+6�/$�b��P   P   7�ӽxE�p���M_��g��{��I5%�VZ��n���}������g���I��� Z��$�����S�^�k|�!��P   P   !���뽢����d��������YF����ϡ�����[��q����0e��ˋ���E��|�g���[d����P   P   k|�V�y��5�d�5ɵ��
�Q_��X��������*��XV��{h��7V�ƾ*��b�������^�����p��[d�P   P   S�^�]�!��"�@�^�氾���WBh��빿.���
h��5�����&���=���g��k�+�����g����g���P   P   �𣾢PW�1�3��kW�C��R���^�Uչ�C�����?x��[�d� ��P�PW��|�����*�����^��|�P   P   ��U��{�T���T��X���DF�4��4s�����]����-0��R��R��)0� {��|���k������E�P   P   �$���Ǿ����i\�B���ĥǾ��$�����p@��`�g�:���0�6�c��cv���c��)0�OW���g��b��ˋ�P   P   � Z����\��q�p�+p��4��U��ѿY�y)����*�yڤ��)�!�Q��Xv��cv��R��P�;��ž*�/e��P   P   �I���y"�ɾų��zKf�Z�����Ⱦ�0"�y
��m6鿀�U�x��ː �!�Q�5�c��R�b� �#����7V���P   P   �g���h=���뾌k���]g�{.g��!��0�꾸�<�%���j��g�x���)��0��-0�[�����{h�p��P   P   ���$M��0����["o�Q�O�2�n�M������,�L�񟢿�j��U�xڤ�:��Z���<x���5���XV�Z��P   P   �}���.M����2W��:nw�PBD�D���v��Ǳ��W�,�L�%��l6���*�^�g���������
h���*����P   P   �n���=��G�Rk��f�z�`H@�9l-���?��-z��Ǳ������<�x
��x)��n@��2s�A��,������̡��P   P   	VZ�е"��뾷P��X�w��o@��&��_&���?���v�M���/�꾄0"�пY�����3��Sչ��빿�X�����P   P   G5%�U���zɾř�&�o�r�D�B�-��&�:l-�D�2�n��!����ȾU����$�BF��^�TBh�O_��YF�P   P   x��GȾrפ�0#���+h�AZP�s�D��o@�aH@�QBD�R�O�{.g�Y����4��åǾ�Q������
����P   P   �g���Γ����$�q��Dg��+h�(�o�Z�w�i�z�<nw�]"o��]g�zKf�*p�A����X��A��氾3ɵ����P   P   �M_��X���U��^]�%�q�1#��ř��P��Tk��3W������k��Ƴ��q�p�i\���T��kW�>�^�3�d���d�P   P   o���"��4���U����tפ��zɾ�뾍G�����0����	ɾ�\������{�T�1�3��"�x�����P   P   xE�|n���"��X��Γ�GȾV��ҵ"��=��.M�&M��h=��y"�����ǾU���PW�]�!�U���P   P   1��zW̽�o��AU��N�����$��R� ف�j����ۛ�����������Q��[�X��aҞ�S�T�]����˽P   P   ��˽̽B���X�Ƽ��31��>�����5᱿�rܿ���e����Aܿ�����x���R>�����J���^X�k�
�P   P   ]�����*���X�G�E�
���U�6����&��W���D��U���D��*���濎Z��!?U�Ĉ
�ے���^X�P   P   S�T��Y��q���T�����?�
��^��{����	�sS��	������읳����D2S�B�	��=��	�]�Ĉ
��J��P   P   `Ҟ�P��A-�I0P�N������qU�ph��Y��Ěx��|���h����
]��Y���]x����=�� ?U����P   P   X��F���P��P�ȼ��f��b>��h����	�[wx�����qh��h>��f>�ka������]x�A�	��Z���R>�P   P   �[���¾(=���7Y��5��e�¾O��n������S�KI��|X�U\O��@a�bO�ka��Y��C2S�����x��P   P   ��Q��@��g]��n�g�m�=������Q��w���������Z?��N>�O8a��@a��f>�	]�����*�����P   P   ������g žՙ��i�e�bx��Q�ľ�S����=�ۿ�sD��M������N>�U\O��h>����ꝳ���D��AܿP   P   ����nb7�p�澈���K�i��xi�_j���L�v�6�~R�����ƆT��M��Y?�{X�oh��h������U�c���P   P   ~ۛ��rF�n+��lި�Ǹt�7LW��Wt��x��������E�Qu������sD�����II�������|���	����D�ޯ��P   P   h����F���������I`Q�&/Q�y\�j�������E�}R��<�ۿ����S�Wwx���x��rS��W��rܿP   P   ف���7�Y��Ř���X���P��@��P�^���j������u�6�����w�������	�W����	��&�2᱿P   P   R�>����d��E���Q��?<�L<��P�y\��x���L��S���Q��n���h��nh���{��4�������P   P   "������ߌžT��'Cu���Q�EA��?<���@�'/Q��Wt�^j��P�ľ��O��b>��qU�~^���U�
�>�P   P   ���Wþ1ء���Agj���W���Q��Q��P�J`Q�8LW��xi�ax��=��c�¾d澲�>�
�D�
�21�P   P   �N���0��շ����n���f�Agj�)Cu�F���X�����ȸt�L�i�i�e�g�m��5��Ǽ��M�������E�ż��P   P   �AU�)�P���P��,Z���n���U��f��ǘ������nި�����ՙ��n��7Y��P�G0P���T���X���X�P   P   �o���� �-���P�ַ��3ء��ž��Y���q+��q��i žg]��(=��P��A-��q��*�B�P   P   yW̽8�����+�P��0��Wþ����@����7��F��rF�pb7����@����¾G���P��Y���̽P   P   r�;������2F�0Γ��ԾC���>�E�j������ҋ�䖅��Cj���>���QԾLS��ZuE��츹�P   P   ��]���e �kI�z>��w�ﾼ�-�q�p�͝����\׿�K׿=������Pp�	T-�.ﾚ̝���H�� �P   P   ��&ٽ�X�EI�������T�A�<0���)ɿ���P$�R�0��7$��t�[�ȿf�rfA�����ڲ����H�P   P   ZuE�`�nz�g�E�)��$��^ I�N]�����i�.�4	o��y��Ko���n��`.��7�g$����H������̝�P   P   LS��t�A�GX!�J�A��{��LT��A��M���b����I�䯚��������Ч��v���+�I����g$��qfA�-�P   P   PԾy�����A���A�񎅾�8Ծ8j-����@W�9�I�!;��Xa����+��4Q��8(��+�I��7�e�T-�P   P   ���W��m�p��J���p��Q�����mp�#�ȿnZ.�|����I����$�.�4���$�4Q��u����`.�Z�ȿOp�P   P   ��>����ێ���_�;�_�}v��*k꾰�>�dy��X�A�n�*���~���4�.�4�*��Χ���n��t����P   P   �Cj���v���+��j�\�����:�������i�u����#��9��y���~���$��� ���Jo���7$�;���P   P   㖅�@z(�C�ؾk���TAh�:h��k���Zؾ�((�V����ֿ�&0��9��)����I��Va�������y��P�0��K׿P   P   �ҋ�c)6�,n�զ��Д|�@*d��=|�M��:�ﾀ�5�Ӏ����ֿ�#�@�n�z���;��ᯚ�1	o��P$��\׿P   P   ����G76��8��4����h�l�\il�D���^&�������5�V��t���X�mZ.�7�I���I�g�.�����P   P   B�j�¡(���𾡫��J틾�{u�H�k��'u����^&��9�ﾷ((���i�cy��!�ȿ=W��b����쿡)ɿ͝�P   P   ��>�G<�9پ�֥������u���m���m��'u�D���M���Zؾ�����>�lp�����M��L]��:0��n�p�P   P   C��7ڸ��x	}��l��,l���m�H�k�]il��=|��k���:��)k꾚��6j-��A�\ I�R�A���-�P   P   �Ծ�ܴ�s������2�h���d��l���u��{u�i�l�A*d�:h����|v���Q���8ԾJT�!�����t��P   P   /Γ�������q�<�`���]�3�h�y	}����K틾�Ҕ|�UAh�k�\�:�_���p������{��(�����x>��P   P   �2F�qB�P�B�v�K�=�`�����󓾬֥�����6���צ��l����+���_��J���A�I�A�f�E�EI�kI�P   P   �������"�P�B���q�t��9ڸ�;پ���8��.n�E�ؾv��܎��n�p���A�FX!�mz��X�e �P   P   
;����ٽ���	qB������ܴ�"�I<�ġ(�I76�e)6�Bz(�������W��y���t�A�`��&ٽ\���P   P   ?K���碽*h��n.�%ā�wԹ������$�y�H�9ic��bm�VHc��cH��N$��e��MM���O���-��l� h��P   P    h��ۦ��N����1�z8��JѾ0�ٻL��#���#�������������-���!bL����S�оrˊ�K1��9�P   P   �l�0%�����i�1�w�����޾t�&�s�o��Ԥ��ֿ:�������/�տ�����Mo� t&� L޾�U��K1�P   P   �-������ ���.�x��>�޾��,�z*��č��,>���/�@�L��L��/�q��M������j�,� L޾qˊ�P   P   �O����)����)�.z��cѾ��&����*oȿ����[��!��{������:~[�Z��9ȿ���� t&�S�оP   P   MM��(�i���)���)��j�m�����to�%k�������m�Kש�x���r���ɩ���m�Y���M���Mo����P   P   �e���
��|�S���2�o�S����i��eL�R���A�&~[��ȩ�I����P��g����ɩ�:~[�q����� bL�P   P   �N$��;����a�I���I��ꅾ��;-7$��僿��տ؞/�����)_���H���P���r������/�-�տ,���P   P   �cH����}����Uo���Q�&o�Ef���^��')H��Ӟ�����XjL�ƚ��)_��H���x��y���ߥL�������P   P   THc���>�ƾ騏�x�n�!�n��v��)Aƾ9����b�[j��}��XjL������ȩ�Iש��!��>�L�������P   P   �bm��, ���޾�料�������!b��x����޾�����l�Zj������מ/�$~[���m��[���/�|:������P   P   7ic�i8 ���羜�������^홾>ٙ�跟�-��4	羬����b��Ӟ���տ@�������*>��ֿ�#��P   P   w�H�S4���޾����D茶����5Q���t��饧�-���޾9��&)H��僿Q���#k��(oȿ���Ԥ��#��P   P   �$�q��_�ƾ�����~���ߴ�AѴ��t��跟�x���(Aƾ�^��-7$�eL�to����y*��q�o�׻L�P   P   �����3ξQ즾�䏾⯌����{d��ߴ�5Q��?ٙ�!b���v��Df����;i�������&���,�s�&�.�P   P   uԹ�(���Pd��F�o��To��E�����~�������^홾���!�n�&o��ꅾ���m��aѾ<�޾��޾JѾP   P   #ā�E�j��T�"hJ�ԧR��To�㯌����E茶��������y�n���Q���I�n�S��j�-z��w��v���x8��P   P   �n.�Us*�{e*�c�3�#hJ�H�o��䏾�����������料ꨏ��Uo�b�I���2���)���)��.�h�1���1�P   P   (h罠������|e*��T�Qd��S즾a�ƾ��޾��羛�޾?�ƾ~�������|�S���)�� �����L��P   P   �碽�㾽����Ws*�G�j�*����3ξs��U4�k8 ��, �������;�
��)�i���)�����/%��ڦ��P   P   �!Z�P(��Fٹ�3��3U�z��/Ѿ����#�:9��@���8�!�#������о_����_T�����븽`]�P   P   `]����nڵ������e��������ڦ%���R�o
z�ψ��ň���y�^R��\%�"3��#2���,e�F�U&��P   P   �븽�u���^�����E1l�����`�pU@�0ဿ�o��M#��p�ǿ�
��H��.����@�h�1����k�F�P   P   ����ƽPFƽ!���e�O��{M�H�O�x�:wſ1���}<��3����`Dſ����O���1����,e�P   P   �_T��/	�)��|X	���T�Ks���G�D�O��w��SUۿfr��7�.ZE�>�6��X�k#ۿO���O�h�"2��P   P   ^���tc?�E4	�i@	�&�?�����e���&@�۫��KDۿ}K�[CT��Gz��@z��1T��7�k#ۿ����@�!3��P   P   ��о�ꂾ��/�=Q�K�/�;�����оke%�㺀�iKſy\�5T��'�������&���1T��X�_Dſ-����\%�P   P   ���0����cf�C1��u1�OHf�s��U���IR�{8���g����6��/z�Q��������@z�=�6����H���]R�P   P    �#�B�׾������d���O�f�d�PД���׾#���y��༿���8E��/z��'���Gz�-ZE��3��
����y�P   P   ��8�y4����vc���t���c��3��g�������8�����Dǿ����6�5T�YCT��7�|<�n�ǿ�ň�P   P   �@��	�frӾT��Uj������@A��0���ӾRM	��~@�����༿�g��x\�|K�dr�.���K#�� ψ�P   P   89�ۚ	���ݾ��о ߾S��%���޾�{о�{ݾRM	��8���y�z8��gKſIDۿQUۿ8wſ�o��l
z�P   P   ��#�(g��ɄӾ��о�c�r�����h��T$�{о�Ӿ���#��IR�⺀�ګ���w��w�.ဿ��R�P   P   ���6ؾ�/��h^���߾̡���%���%�h����޾0��g�����׾U��je%��&@�B�O�F�O�nU@�ئ%�P   P   ,Ѿ%鬾�9��4����l����������%����%��@A��3��PД�s����о�e���G�yM��`����P   P   x��!T��wg� [e�<����������̡�r��S�𾧨���c��f�d�NHf�:������Js��M���������P   P   �3U��2@��0�92�3jP�<����l���߾�c�߾Vj���t����O��u1�K�/�$�?���T��e�C1l���e�P   P   3�h�	�t�	���:2�"[e�4���i^����о��оT��vc����d�C1�>Q�i@	�{X	� ��������P   P   Eٹ��.ǽ���u�	��0�yg��9���/��ʄӾ��ݾgrӾ �������cf���/�E4	�)��OFƽ�^��lڵ�P   P   P(��q(���.ǽi�	��2@�"T��'鬾�6ؾ*g��ݚ	��	�{4��D�׾1����ꂾtc?��/	��ƽ�u�����P   P   -���$�h̀��н!!�s�k����gԾA�i��n5�d��i� �M�Ӿ�����k�!f ���νG��� $�P   P   � $��p$��|��7׽�m/�C����g���W���� ���<��`M��SM���<�ِ ����������.��*ֽ�8{�P   P   G���7G��^��0�ֽ��4�뎾�sӾ�M�i�A���n��B�������2��Tn��RA����Ҿ7����F4��*ֽP   P   ��ν�����.��riϽ�2/�Jڎ��4۾���q.Z�ԇ���/��K���U�������e����Y������ھ7����.�P   P   !f �2lƽ�z��N�ƽ�� ��T��hMӾ���}Ic�ᚿt�ƿ���f��^��Ĳƿ#����c�����Ҿ���P   P   �k�E�>ɽ8Vɽ�j�`_k�?"��,�Z��ך��uѿ4��(��O��e��9]ѿ#�����Y����P   P   ����wM�?
�s���C
��-M�k�������)aA�9n��C�ƿ�������*����d��Ĳƿ�e���RA�����P   P   L�Ӿ�	���D��l��b��D�����Ӿ�� ��Fn�\����z���*���*�N��]�����Tn�ؐ �P   P   h� �Ⱥ��.鉾@1n�xd���m�0���ǆ���� ���<����du������y����'��e��T����2����<�P   P   c���ؾ�+�����{���ݐ���䯾N޵���ؾ��M�����du�������3�����J��������SM�P   P   m5�Q����ھ�}�}6	��A��	�$��gھI���M����\��B�ƿ�uѿr�ƿ�/���B���`M�P   P   g������G�N���r7�9Z�u)Z�xJ7��h�	��I�����<��Fn�8n���ך�ᚿ҇��~�n���<�P   P   @��پ��ھ.���'K��ć�"�������K��h��gھ��ؾ�� ��� �(aA�Z�{Ic�o.Z�g�A��� �P   P   eԾSR4���^��W7������Ʃ�ǩ�����xJ7�$�M޵�Ɔ���Ӿ����,��������M��W��P   P   ����Q���	������	�Z�#���Ʃ�"��u)Z��	��䯾0������j���="��gMӾ�4۾�sӾ�g��P   P   p�k��M��1E�XVn�����1'�Z������ć�9Z��A�ݐ����m��D��-M�^_k��T��Iڎ�뎾B���P   P   !!����
����̤d������	��W7��'K��r7�}6	�{���xd��b��C
��j��� ��2/���4��m/�P   P   �нحǽ�tʽ�����YVn�����^�.��O���}����A1n��l�t��8VɽN�ƽpiϽ.�ֽ�7׽P   P   g̀�Q���+����tʽ�
��1E��	��S4����ھ�G���ھ�+��/鉾�D�?
�>ɽ�z���.���^���|�P   P   ��$��|H�R���ڭǽ	���M��Q��U�پ���R���ؾɺ���	��xM�E�3lƽ�����7G��p$�P   P   �|�L�n�9'�j+~��ؽB�'�Orp�=���SǾ ��N�㾲�ƾF����o��'�J]׽|������k�P   P   ��k�?Jm�E| �o煽|�e>�ۅ��')����뾿(
�������Q
����κ�&��C�=��C��������P   P   ���Mj��;i�@��������?M��9����־I��p�)���?�N�G���?�_�)�g���q־9֙�#�L��������P   P   |�9�Ў�}���$M��+��(��x��9�F�I�j������|j�fF�il�1��џ�"�L��C�P   P   I]׽$�n���/� To�-�׽M>�l��#��^�"��|W��p������\��r옿:]���NW��"�1�9֙�B�=�P   P   �'�`ý0���󚀽'�ý�M'�^Q��9�־L���qW��v���������������Lf���NW�il��q־&��P   P   ��o�ڋ��Lѽ&'��rPѽ�����o��㺾���vF�e����yOÿ��ͿLÿ���9]��fF�f��κ�P   P   F����`�B5.�&%���.�W�`�7��\v��)�wj��蘿�����Ϳ��Ϳ���q옿~|j�^�)����P   P   ��ƾD|��O���x����������N��KE��l�ƾ��	�Ԩ?����O������yOÿ����\��~����?�P
�P   P   ��㾐���l�Ⱦ���4��#��7��EȾ,����E�<����G����蘿������������M�G����P   P   N�ڡھ�C���.��fc�tx{�7c�?�-������1ھ���<��Ө?�wj�e���v���p��G�j���?����P   P   ���3�ھ5�
���V�PB���q˿�b˿���zV�F�
��1ھ�E㾧�	��)��vF��qW��|W�7�F�n�)��(
�P   P   QǾ<����#����V�C����Up��������zV�����,���l�ƾ\v���K��]�"�w��G�����P   P   <���`���9�Ⱦf�-�`!�������(�W�(�������?�-��EȾKE��7���㺾8�־!��&����־&)��P   P   Mrp�`Qa�<z���8��c�$D˿d���(�Up��b˿7c��7�N��V�`���o�^Q��j���+���9��څ��P   P   @�'�
�@g.�o���K ��*{�$D˿������q˿sx{��#�����.�����M'�L>��$M��?M�	e>�P   P   �ؽ�{Ľ�ҽTF��{��K ��c�`!��B��OB���fc��4�������rPѽ'�ý,�׽｡���|�P   P   g+~���p��y���߳�TF�o����8�f�-���V���V��.���w��'%�''��󚀽 To�}�>���n煽P   P   7'����2�1��y���ҽAg.�<z��9�Ⱦ�#��5�
��C��l�ȾO���C5.��Lѽ1�����/�Ў�:i�D| �P   P   J�n���������p��{Ľ
�aQa�`���=���4�ھڡھ����E|����`�ۋ�	`ý'�n�9�Mj��=Jm�P   P   &��<�`@<U⠺kļ��l��fս�'���l�b���Is���v���k��/똾<sl��&��eԽ��j��z��B�n�C<P   P   C<��A<%�~��ۼ�������$:�+�������dľN�վ��վ�Bľ楾�c���9��a𽱯���׼T/>�P   P   �n����;B��\wڼ��������P�x����+��3�&������W�������m��NcO��:�����׼P   P   �z����4�Xb9�G¼�j��[��K�X�񜟾��׾k���>�15+��,+�g'�)n�l�׾�K��=X��:�����P   P   ��j�����dN)�o���4�k����O�����z��l���52��I��fQ���H��2�=t��9��K��McO��a�P   P   �eԽhz_�q���������_���Խ=�9�ܝ����׾�����9��mZ�K�m�_�m�6]Z��{9�=t�k�׾�m���9�P   P   �&�7ٽO��r(��j��"ٽλ&��u�������}�+)2�ChZ��w��r��-�w�5]Z��2�)n������c��P   P   ;sl��8�Ŏ%��#���#�oX%���7�Pl��ߥ�/�龌(��H��m�hr���r��_�m���H�g'�V��楾P   P   /똾�'���ʗ�V��]���䮾<����⊾f����ľ���� +��\Q��m��w�K�m��fQ��,+����BľP   P   �k��n(��"���$�)�G��G�Z�$�/U�N���?��߇վ���� +��H�BhZ��mZ��I�05+�����վP   P   �v���ؾ�u"���춿�oο����ȁ�
"��*ؾ���߇վ����(�*)2���9��52��>�&��M�վP   P   Hs����ؾ�$4��P���	��,�ԣ,���<����3��*ؾ?���ľ.�龩}����k��j�� 3꾯dľP   P   a�������P"�G;���f��`��Q��ܸ`��L�<��
"�N���f����ߥ�������׾y�ྶ�׾�+�����P   P   ��l������1ҁ������`�+s���r��۸`���ȁ�.U�⊾Pl��u��ܝ������𜟾w���*���P   P   �'�%,8�c���m$�_����,��H��*s���Q��ԣ,�����Y�$�<�����7�λ&�<�9��O�I�X��P�$:�P   P   �fս��ٽEz%����asG��(ο�,���`��`��,�oο�G� 䮾oX%�"ٽ��Խ��Z��������P   P   ��l�� a�x���p#��0��asG�_�������f��	�춿(�G�]�����#�j����_�4�k��j����������P   P   gļ��I� �ހ���p#����m$�1ҁ�G;���P������$�U���#�s(������r���G¼Zwڼ�ۼP   P   :⠺��K��/�I� �x��Ez%�c�����P"��$4��u"�"���ʗ�Ŏ%�P��w���nN)�nb9�G����~�P   P   �`@<Q��;�K���� a���ٽ&,8���������ؾ�ؾn(���'���8�9ٽlz_������4����;��A<P   P   %�=܍=��<�<j����_�bؽ��+�sn��I��or��EN��.n�2�+�e�׽kV^��9����$<�F�<�=P   P   �=��=��<G��;#���^�v�Z޽�K'��`��ᇾ:���Ҷ���̇�-�_���&��yݽ� u�0�����<1q�<P   P   �F�<n�=H�<��;@�¼X/���W����;��|�����uӮ�����������f�{� $;�7K���=��ƿ���<P   P   ��$<y��<o�<�{!<V�������4�K��׌�T�����Ͼ�<��0�C�Ͼlɱ�_���{"K�oN��=��-���P   P   �9��Ib<���<?�<<݆�c<v�\����K�]�������|8� ����%����m^���z��{"K�6K��� u�P   P   hV^����[����B������e�^���ݽ�u;��ǌ�����ɵ򾦘�� �a����|��m^��^��� $;��yݽP   P   d�׽@���
�p���b��p��͔�j�׽�'���{��屾�*�*��2?�	�%��9�����lɱ�f�{���&�P   P   2�+��&���&�-�5���5�Y�&����s+��_�4���N�Ͼ�������%��%�a��%��C�Ͼ����,�_�P   P   .n��%��H%����ھ��b|ھ����]̃�A�m�c��������&������2?�� � ���0�����̇�P   P   EN�����������[���������[�2h�p������{����ﵾ�&����*����� ���<����Ҷ��P   P   pr��q��~M��)�����Մ�߰��ϳ���L�7�����{�������N�Ͼ�*�ȵ�{8龽�ϾuӮ�:���P   P   �I���[�^f��c迻LA��l{��U{�~A���)�e�7������c���4����屾��������S�������ᇾP   P   sn�t��:EM��D��\�Ϣ�{���¿��*X\�����L�o��A�m��_���{��ǌ�]����׌��|��`�P   P   ��+�����p���⳿2%A�Ţ�B���@��¿��}A��ϳ�2h�]̃� s+��'��u;���K�3�K���;��K'�P   P   bؽ�	��ë��s[�ĝ�/;{�^���B��{����U{�ް���[��������j�׽��ݽ[������W��Z޽P   P   ��_��'��g�&��1ھgƉ�5V�/;{�Ţ�Ϣ��l{�Ԅ�����a|ھY�&��͔�f�^�c<v���W/��\�v�P   P   j���T��y�p���5���gƉ�ĝ�1%A���\��LA����������5��p�����?݆�W��?�¼!���P   P   �<�1<�i����b���5��1ھ�s[��⳿�D迈c��)����[���ھ,�5���b��B��4�<�{!<��;J��;P   P   ��<ϡ�<ly�<�i��x�p�f�&��ë�p��9EM�^f��~M����G%����&��p�w���< o�<E�<��<P   P   ܍=��=ϡ�<�1<�T���'���	�����t���[�q⾅����%���&�A������;b<t��<l�=��=P   P   	�n=�e=�3J=p?=�~�<x���|�|�h�����;�\Tp�U���Kop�q�;�����|����[߃<`=�K=�Gf=P   P   �Gf=�
f=��J=Wc=1%n<.p�٬S�H½��v�6���M�4�M��n6����K����lR��Pj���s<�z=7K=P   P   �K=�b]=L�J=l�=��T<�b��U1m�x�ѽi���@�8�]�9/h�&�]�3�@�h�p�н�~k��V��uZ<�z=P   P   `=�7D=�D=L�=�wo<���k|��`�U/)��7\��*��d?���6�����}�[���(�b����z��V����s<P   P   a߃<
=�`!=��	=Ǐ�<�^n�^�l��I�{�0�IKo�D���B(����,��=����n�X�0�b�併~k��Pj�P   P   �����;��c<��c<k��;�[���S��sѽ�)�!Ao������@�����f����+���Ԙ��n���(�o�н�lR�P   P   �|�ZkC��*<���?�3�;��C�,|�+����=��\������>��C�ɾ�Ѿ=�ɾ�+��=���}�[�g�K���P   P   �����]�(���D���D�In(����7��y��8�@�����!��I�����Ѿ�Ѿf���,�����3�@����P   P   r�;��:~��Ȼ����L��-f��M���a}�D);��-6�l�]�13������I���C�ɾ������6��&�]��n6�P   P   Mop��¾���&��Â�D覿�ʦ����� W&������o��gM���g�13���!���>���@��B(��d?��9/h�5�M�P   P   V���rA�,�m�҅ٿ1t�?u5�bI��ٿ�m�j{龊!���gM�l�]������������D����*��9�]���M�P   P   ^Tp��$����u���l�X��`I��09l�
p�M���j{龶�o��-6�8�@��\� Ao�IKo��7\���@�v�6�P   P   ;������tm�ۢ�׆�f��/���V������
p��m����D);�y���=��)�{�0�T/)�i���P   P   i����}��|&��2ٿ�Sl��^���}��|���V��09l��ٿW&��a}��7��,����sѽ�I彟`�x�ѽ�H½P   P   ~�|��@��J��u��:��?��-���}��/��_I��aI�����M����.|��S�_�l��k|�U1m�ڬS�P   P   {����pC��M(�,��*����C5��?���^��f��X��>u5��ʦ�,f��In(��C��[���^n����b��!.p�P   P   �~�<̙;]�;�CTD�Ee�*���:��Sl�׆��l�0t�C覿K����D�5�;�O��;���<�wo<��T</%n<P   P   o?=k'	=�b<�<?�CTD�+��u���2ٿڢ�t��хٿ�Â������D�·?���c<��	=I�=j�=Wc=P   P   �3J=jUC=�� =�b<\�;��M(��J���|&�~tm����*�m���&��Ȼ�\�(��*<���c<�`!=�D=J�J=��J=P   P   �e=��\=jUC=k'	=̙;�pC��@��}������$�qA��¾��:~���[kC���;
=�7D=�b]=�
f=P   P   z��=A��=���=�/e=;�=js<<���Bު����|_E��_Y��E����0��#C�_�><�| =�f=�׆=���=P   P   ���=@��=��=U�e=�<&=C�<"�(���8�%i��4+�:�	��	��뽜2��V8�0�%��9�<�I'=ܥf=�;�=P   P   �׆=�?�=���=z�e=�#=�v�<�4�WG2��ɝ�#N۽�L�I��8���ڽ�Y���1��q/�tܐ<��$=ݥf=P   P   �f=Ms�=�]�=J�e=v&=Z��<JZS�?eF�*믽�c����p�&�E�&�nx�����dK���E���N�vܐ<�I'=P   P   �| =��O=�x^=&QO=��=���<�3�OGF�LY����y},�pE��<N��TE��J,��]�Ÿ��E��q/��9�<P   P   f�><��<u3�<:.�<�ȼ<<�=<e'�I�1�tί�Û���4��X��vk�jk���W�{�4��]�dK���1�-�%�P   P   $C𼞭�:��Yh��H���較��M/8������<��^u,��X�Y)v�Bp���v���W��J,������Y��V8�P   P   2��(�.Q!��C�H�C�s� �r=�p������� ۽���EkE�{k�Os��Bp��jk��TE�nx���ڽ�2��P   P   �����j�������� ��{��}j��X����!�^�&�gBN�{k�Y)v��vk��<N�F�&��8���P   P   �E��̵�
x(�D������.�����'�����D��*	���
�^�&�EkE��X��X�pE�q�&�J��	�P   P   �_Y����Gq���߿�8$�w�:�v	$��߿؁p����X��*	��!����^u,���4�z},����L�<�	�P   P   ~_E���ᾫE��+��sas�~�������s�&H��ㇿ���D���� ۽�<��Û����c��%N۽7+�P   P   �������q�Q��˯�������T��e���K���&H�ׁp�����X���������uί�MY��+믽�ɝ�(i��P   P   Eު��_j��(��:߿�8s�4���O%���!��e����s��߿��'�|j�p��P/8�K�1�PGF�AeF�ZG2���8�P   P   ����q��~��r����$����hT��O%���T�����u	$�-����{��r=潉��"e'� �3�RZS��4�/�(�P   P   ^s<<�鼎� �� �������:����4�������~���v�:��
� �r� ����,�=<���<U��<�v�<>�<P   P   9�=sT�<����VC��7������$��8s�ʯ��ras��8$������G�C��H��ȼ<��=v&=�#=�<&=P   P   �/e=��N=]��<J���VC�� �q����:߿P��*����߿D����}�C�Zh�2.�<!QO=F�e=w�e=S�e=P   P   ���=� �=�^=_��<����� ��~���(� q��E��Gq�	x(����-Q!�:��o3�<�x^=~]�=���=��=P   P   @��=��=� �=��N=xT�<���q��_j������������̵���j�(罞�鼙�<܎O=Ks�=�?�=?��=P   P   r��=t�=�ƙ=Vۉ=B�Y=ŀ�<v`ܻ[�`�j�ݽ	�t�-��,��0޽;a�w=ܻ�!�<�$Z=�(�=��=���=P   P   ���=���=��=`9�=CSi=�$=u�<[F7�^	,����ܯ�y߯�����+�)�5���<��$=�j=S��=��=P   P   ��=�h�=ߙ=0C�=<j=�=(=G�<�l�"��ucS��݊��施Ê��R�_��s_�m@�<{')={k=T��=P   P   �(�=�g�=3W�=6��=�vi=9P(=ף<W<��X��g��e���O���;��q)���`f�Qe �E�����<{')=�j=P   P   �$Z=�v=�=��v=q�Y=7=$=���<\����K�<-��yC����ֽ��⽜�ֽ!󳽄���_
�E��n@�<��$=P   P   �!�<W7==�=�6=k��<���<9?i��1�(&���Ҿ��｣��g������z������Qe �z_���<P   P   �=ܻ?�\��ü�Y�1¼�qZ��ٻ��5�"���f�B:��0�o���7�������"󳽬`f�c��0�5�P   P   @a�f�����n/�tE/���������_�>W+���R��J��4�ֽy��7=��7�g����ֽr)��"�R�#�+�P   P   �0޽y�I�а��_���O���澟3��=�H��ݽ\��������=��+��y��p�������⽥;��Ê����P   P   �,�*f���&�cm��#����o�l���������q�S3�������=��4�ֽ1��ｬ�ֽ�O���施}߯�P   P   x�-��Xžt�T��)ÿ����"�l����¿Y�S���ľ�-�S3�������J��C:���Ҿ�zC���e���݊��ܯ�P   P   �	�?ž�qo�����+�R����|���XR��A��H�n���ľ�q�]�����R���f�)&��=-���g�zcS���P   P   o�ݽ�)��kQT����BJp��[��>����B����o��A��X�S������ݽAW+�"뼈1��K�X�-��f	,�P   P   c�`�I����¿=�R�BV���/��X+���B��WR���¿���=�H���_���5�n?i�t���q<��U�l�sF7�P   P   �`ܻR���6?��ɔl����'���о���/��=���{���k��n�l��3������.�ٻ���<���<ף<	G�<u�<P   P   ���<r{Z�Ä�[_�E䖿�e"�'���AV���[�����߁"���������qZ�b��<2=$=6P(=�=(=�$=P   P   ?�Y=j'=P����.�s�D䖿���<�R�AJp�)�R�����#���O�sE/�1¼�6=l�Y=�vi=	<j=@Si=P   P   Uۉ=��v=G(=�輏�.�Z_�Ȕl��¿��������)ÿam�\���n/��Y��=��v=4��=.C�=^9�=P   P   �ƙ=+0�=Ę=H(=P���5?����iQT��qo�r�T��&�ΰ�����ü=�=1W�=ߙ=��=P   P   t�=�?�=+0�=��v=m'=_{Z�O���I��)��?ž�Xž(f��v�I� f��:�\�U7=�v=�g�=�h�=���=P   P   �l�=���=EC�=�ӑ=��q=ny=${�;��	��ՠ�ή�>��G��p*��]5
�MC�;
�=�	r=��=�o�=宥=P   P   宥=
��=ƪ�=���=���=�[Q=}�=ϟ<͊�����JoU�zU����Ax���X<F�=��Q=K;�=84�=�Ѡ=P   P   �o�=�e�=FR�=���=�Ʌ=-\=&�=���<��:5\��ڢ���	��^�dυ�N!�:<�<��=4�\= �=94�=P   P   ��=���=��=��=���=$7\=%� =Y�<�g+;�V{�p��7��@������0y��q6;Q��<�W!=5�\=L;�=P   P   �	r=��=�q�=#�=��q=bqQ=i�=��<���:�w��й��C��%T���B�	=��-��7d;Q��<��=��Q=P   P   �=K�!=�C=.K=A "=��=w�=���<c-;�g����\ga��ꂽKڂ��a�ؔ��-���q6;;�<F�=P   P   =C�;��3��f�o���
e��p+��4�;��<�:�z�����ka�b��nF���F���a�
=��0y�!�:�X<P   P   b5
��f�����_�B���I�Y���_$	��l������(\�	#C�+����O��nF��Kڂ���B����lυ�Jx��P   P   t*���� �Eņ�)h��Euξ���^�����m5�� ��#������AT�+���b���ꂽ�%T�D���^����P   P   M�뽜�}�7���8���g��g�n�7�����u|�'�꽲KT��+	����
#C��ka�^ga��C�<����	�zU�P   P   A������Ly%�,l��0)տ�����Կ>����$�%�����KT�%��+\񼴮���Թ�y����SoU�P   P   Ԯ�����w9��O��k����H��H��e�q޻���8�%�'��"������)�z��g���w���V{�B\�����P   P   �ՠ�S*}�nQ%��=��&�0��_��ԅ���H��Kx0�q޻���$��u|�n5���l����:1-;}��:Eg+;��:݊��P   P   ��	��" �31�LB����R\��LΨ�=ƨ��H���e�=����꾏��a$	���<���<��<Q�<���<��<P   P   �z�;ǎ��m��[�7���Կ��H�����LΨ�Ӆ��
�H���Կm�7�^��Y����4�;s�=e�=!� ="�=w�=P   P   iy=��*�|�0���9fg�cv���H�R\���_����H����g�����I��p+���=]qQ= 7\= -\=~[Q=P   P   ��q=�"=DQc����ξ9fg���Կ��%�0�i��/)տ��g�CuξB���
e�= "=��q=���=�Ʌ=���=P   P   �ӑ=��={=>���/���Z�7�KB���=���O��+l���8�'h��]�o��*K=!�=��=���=���=P   P   DC�=�m�=�e�={=9Qc�y��m��21�lQ%��w9�Jy%�4��Cņ�����f��C=�q�=��=ER�=Ū�=P   P   ���=dK�=�m�=��=�"=W�*�]̌��" �P*}����������}��� ��f��m�3�I�!=��=���=�e�=	��=P   P   Ɵ=f�=we�=~O�=�1l=�"=ȋW<����?k��4��yJȽ�e����k�����Z�V<t�"=LYl=_l�=`��=�)�=P   P   �)�= �=�U�=A��=���=fZ=h�=��<�\��먼X��a��3$���q��
�<�=�Z==�$�=�o�=P   P   `��=��=�l�=���=��=�(j=�;=��=���<z�5;�?���1����Ve8;J$�<�U=��;=]�j=z��=�$�=P   P   `l�=�b�=[�=�R�=���=e,j=_7A=�!=t��<���;�]5�%�³���1�0m <
��<`�=��A=^�j=ﷃ=P   P   MYl=��s=)�u=a�s=U0l=kZ=1#;=2(=�ͮ<�7�;����V�X�/����0X�ʨ��"��;Xٯ<`�=��;=�Z=P   P   t�"=6$=)S=�\=�6=	�"=��={=Y��<�^�;��λ��R���ӿ��z����˻��;��<�U=�=P   P   R�V<=�;����X�L�;Q;
X<�\�<��<���;�T��p��?�׼��|C׼�z��ר��'m <E$�<�
�<P   P   ������V���`�W)ὔ����gU��ڪ��]�U`:;	t3���X��,���5���ӿ��0X��1�e8;=r�P   P   ��k�����%P�vR���t��
��{�O�̽��p@j�����,�ߥ��ބ��,��A�׼V��4���ӳ���A$��P   P   �e���)C�5Ű�6���$��f$���p:���WB�f��� ��U0�����X�s����c�X�8���1�i��P   P   JȽ��p��;�uM�uԏ��o��<���z�L�<}�L�o�=Hǽ� ��,�!t3�U����λ�����]5��?�a��P   P   �4����p����3n����̿���:��\�̿�$��-��L�o�f�����2`:;��;�^�;t7�;y��;�5;�먼P   P   �?k��B�S	�c���n���'��o>���'����$��<}�WB�q@j��]���<S��<�ͮ<k��<���<�\�P   P   ����;���}��6CM�g�̿g�'��`X��TX���'�\�̿y�L�o:��̽���ڪ�|\�<x=/(=�!=��=��<P   P   ��W<��U��O����ն��^���v>��`X��o>�9��;�����z�O��gU��	X<��=-#;=[7A=�;=c�=P   P   �"=�;�\������R$��`��^��g�'���'�����o���f$�	������Q;�"=kZ=a,j=�(j=fZ=P   P   }1l=X=���3��:���R$�ն��f�̿�n翣�̿tԏ� �$��t��V)�"L��6=P0l=���=��=���=P   P   }O�=:�s=��=iV�2�ླྀ�����5CM��c��2n���uM�4��tR��`��X��\=]�s=�R�=���=?��=P   P   ve�=�S�=��u=��=����\���O��}��Q	�����;�3Ű�%P������'S=&�u=[�=�l�=�U�=P   P   f�=�q�=�S�=<�s=X=�;��U��;���B���p���p��)C�������V�T�;5$=��s=�b�=��= �=P   P   ���=�ތ=FC�=�Rw=��M=�=�d2<鸓��E�&����<��Q뒽��E�J����1<zf=@�M=lhw=�P�=��=P   P   ��=k��=r��=㷂=9�l=7(F=N=�Q�<y/�:
�m�O"¼G¼�Mn��z:,�<�=AIF=��l=�΂=�Ή=P   P   �P�=ᯈ=�D�=ض�=Êt=��Y=�4=�=c��<<���:&\庎��:W<x7�<�5=�5=�0Z=I�t=�΂=P   P   mhw=��{=x�{=�Hw=��l=t�Y=��==��=���<N�<�#<&՚;�:�;Ʋ<�<^�<O=��==�0Z=��l=P   P   A�M=L�O=��O=ҶO=��M=!F=��4=��=���<�!�<_�(<�k�;08;ol�;��)<(Û<}C�<O=�5=AIF=P   P   zf=�r�<���<!�<̤�<�y=�=;=���<�)�<�$<y1;%(��η���4;��%<&Û<^�<�5=�=P   P   �1<	S
�T'.�Jp�B�,�yLݹ!�2<���<�<�<�w�<��(<�a1;6�C���t�A�|�4;��)<�<s7�<,�<P   P   R���[�;�̿��<羽}���WR��E�:�j����:<2�<u�;k����p����Bη�^l�;��<�V<�z:P   P   �E��Ͻ��(��`���v�N`��>(�Z"νW\D��\k�z�:r��;��;w���D�C�X(��8;�:�;�:�Mn�P   P   U뒽�.�����"ɾ���z��Ⱦ뺉���i��ɒ��ƨٺn��; u�;�a1;�x1;�k�;՚;�\�+G¼P   P   �<����@���+���I�<(`� vI�]�䈷�@��p��ʒ���y�:-�<��(<�$<R�(<�#<佢:_"¼P   P   +���U�@��uʾ�5�u�������F��V�5���ɾ@�j���\k��<�w�<�)�<�!�<N�<�<'�m�P   P   �E�S��跾��5������(߿�i��߿ʛ�V�5�㈷���X\D�g�:�<�<���<��<���<X��<�.�:P   P   �����|ν�艾>���e��r"߿3b�[�߿�F��]�뺉�Z"νn��}��<8=��=��=�=�Q�<P   P   �d2<�:��M(���Ⱦ�I������n��3b��i��� vI��Ⱦ�>(�G�:��2<�=��4=��==�4=I=P   P   ��=*,ȹ(���(`��[�`�����q"߿�(߿���;(`��z�N`�WR���Mݹ�y=!F=q�Y=��Y=3(F=P   P   ��M=L =�9+�;P����v��[��I��e������u��߬I�����v�|���I�,�Ť�<��M=��l=��t=6�l=P   P   �Rw=��O=ű�<�{m�:P���(`���Ⱦ=����5��5�*���"ɾ�`�;羽Lp��<϶O=�Hw=׶�=ⷂ=P   P   EC�=��{=p�O=Ǳ�<�9+�(���M(��艾跾�uʾ�������(�ʿ��R'.����<��O=u�{=�D�=r��=P   P   �ތ=���=��{=��O=N =#*ȹ��:��|νQ��S�@���@��.��ϽW�;��R
��r�<J�O=��{=ை=j��=P   P   z�k=oAh=�\=�E=R�=���<ҹ�:��ǼLQP��������A��b�P�B�ȼ���:��<]~=�E=��\=;Fh=P   P   <Fh=/@h=n�b=}�U=�4?=�=�J�<ͯ7<ʖ�+���Jؼ�xؼk~�������6<��<]�=jA?=%�U=Ϭb=P   P   ��\=��^=;�\=��U=��H=j#3=�h=Cd�<�!�<0,�;�"��Y�?��f�����;��<�x�<@=�@3=`�H=%�U=P   P   �E=/G=�)G=|	E=�(?=�3=�y=�=���<+f�<��,<Ɂ�;^��;�
-<*��<��<x�=�=�@3=kA?=P   P   ]~=xF=w�=�H=�=��=�e=�=���<��<�bg<� <�&<� <R�g<��<,6�<x�=@=^�=P   P   ��<=i�< �<�8�<���<fN�<�A�<}q�<p��<厥<�s<2�%<*�;i�;�&<?�s<��<��<�x�<��<P   P   ���:pW)�����tż���+�'�8�:'	8<�Z�<���<>�g<R�%<{�;gɶ;��;�&<M�g<&��<��<��6<P   P   I�ȼ�GO�񙜽�4��)���9���aN��Ǽ�������;�E-<N� <���;���;dɶ;i�;�� <
-<���;����P   P   h�P���ɽ�
��[L��_�DL�_����Ƚ*�O����f�� ��;�1<���;{�; �;�&<D��;�h��u~��P   P   �A���Q�{#w�R!��.�ӾljӾ�د��v�e��������ּ}�9���;L� <N�%<,�%<� <���;��?��xؼP   P   ���C~0��͡��6 �;�,��*@�]�,������d���/��h����ּ����E-<9�g<�s<�bg<��,<6%���JؼP   P   ���lh0�g���3�]�q��*�����&�q�q�������/�����������;���<Ꭵ<��<$f�<,�;7��P   P   RQP�-�Ȭ���%�k�����˿T�˿����q���d��e��,�O������Z�<l��<���<���<�!�<=ʖ�P   P   ��Ǽ�
ɽݿv�� ���q���˿m�<g���˿%�q������v���ȽǼ	8<xq�<�=�=;d�<��7<P   P   I��:�aN���ܯ��,����	�m�T����]�,��د�_���aN���:�A�<�e=�y=�h=�J�<P   P   ���<D�&�����K��CӾb
@�����˿��˿�*���*@�kjӾDL��9��4�'�aN�<��=�3=h#3=�=P   P   P�=�2�<q�������^��CӾ�,���q�k���]�q�;�,�-�Ӿ�_�)��������<�=�(?=��H=�4?=P   P   �E=7y=���<�ü�����K�ܯ�� ��%��3�6 �Q!���[L��4��uż�8�<�H=z	E=��U={�U=P   P   �\=�BG=2=���<n�������ܿv�Ǭ��f���͡�y#w��
�𙜽�����<u�=�)G=9�\=m�b=P   P   nAh=˓^=�BG=9y=�2�<7�&��aN��
ɽ,�jh0�A~0��Q���ɽ�GO�lW)�<i�<vF=/G=��^=.@h=P   P   4@0=�|,=��=�=zG�<��<b�N� �"��{�������|����?������
Q��	<�Ҽ<��=��=^x,=P   P   ^x,=x,=^'=ٟ=�=���<ۍO<Q������n�4��L���������N<IN�< �=ۚ=)'=P   P   ��=��!=D�=1�=٢=�W�<{��<�<�[�;���!���5����т!��n�;�S<r�<yQ�<�=ܚ=P   P   ��=#=n=
�=�=-K�< }�<�ʵ<��<�|!<���;(�:�!�:Q��;�!<��<Wյ<\��<yQ�< �=P   P   �Ҽ<J��<JG�<�в<���<�l�<�~�<N͵<R�<�m<��&<\l�;:��;���;'<�Mm<�*�<Wյ<r�<IN�<P   P   �	<eB;�'�-��CE;v�<edO<��<��<�#m<L�><R;<u�;v��;�s<`�><�Mm<��<�S<��N<P   P   �
Q�;м����y!��H��&ϼK,O�ob���5�;��!<G'<0K<tv�;��;��;�s<'<�!<�n�;���P   P   �����������J׽�$׽�S��M��n��3���"8�m�;��;��;���;��;q��;���;C��;��!�����P   P   �?����߽"1&���S��f�t�S�)�%��޽a[�Bq�,����:�S�;��;qv�;u�;/��;c!�:�����P   P   ���`����|��u��k־�L־9-��T8|��y���������3����:��;.K<N;<Ol�;��:�5��L�P   P   ����S�7����w���5�(yL���4�[^�ʌ��?B7�_������,�h�;D'<H�><��&<���;/��4�P   P   ~����7��:���R!�Є�{5�������!��ֲ�?B7����Dq�28���!<�#m<�m<�|!<���
n�P   P   &��>���У�6A!�tؘ�L� ����q �����!�ʌ���y�b[�6����5�;��<O�<��<�[�;���P   P   $��߽Bn|��w�����&� ��UG��JG�q ����Z^�S8|��޽o���b����<J͵<�ʵ<׬<����P   P   n�N�PE���%�*��4�4����&���UG��������4�9-��)�%�	M��R,O�]dO<�~�<}�<w��<ЍO<P   P   ��<��μ��E{S��־HKL����&� �K� �{5��'yL��L־t�S��S���&ϼn�<�l�<)K�<�W�<���<P   P   wG�<cJ;L����ֽ��e��־4�4�����tؘ�Є��5�k־�f��$׽�H�fCE;���<�=آ=�=P   P   �=I�<�H�*� ��ֽD{S�*���w�6A!��R!�w���u����S�J׽�y!����в<�=0�=؟=P   P   ��=C;=�ܮ<�F�K�����%�An|��У��:�������|�!1&���������'�GG�<l=B�=]'=P   P   �|,=X�!=C;=I�<{J;��μOE���߽=���7�R�7�_����߽����9мeB;H��<"=��!=x,=P   P   � �<���<�l�<
��<�Z�;����(LZ�f��9$ƽa�Խ�Uƽ������Z����������;7M�<�8�<���<P   P   ���<���<���<��<1��<_�<��;��ֆ�	���Z1��O��'O�h1�@W��R�����@�M�<�E�<��<B��<P   P   �8�<b�<MD�<9�<���<��z<͢<��:r�㻴�v��W��� ������Hw���廨��:�<�3z<l�<��<P   P   8M�<���<���<�g�<,m�<��z<U`R<��<�ʃ;1�����s�����􆸻���p�;z<R<�3z<�E�<P   P   ���;�͚;נ�;�q�;���;�z<=�<�<���;�U�;��:��s�t�kus��e�:,�;�k�;z<�<N�<P   P   ��� >k�����g���Zj�����<�)��:,�;ؐ�;*�[;f��:��r:
�r:���:î[;*�;m�;���:��@�P   P   ����L.��1Y��vi���X���-���U������Ù��!�:���:FR�:d3�:6�:���:�e�:(������T���P   P   ��Z����� ٽ���F}����ؽ�2���Z�{
��2�u�a���E@m�|u:Yn�:a3�:��r:�us������Hw�DW��P   P   ����������6���d�7�v��Id�<(6�>7����i�0�혪�������|u:AR�:��r:��������h1�P   P   �Uƽ,�+�����O0�����H���⻾d��"+���Ž'PN�������P@m����:W��:͝s�y��� ���'O�P   P   c�Խ�KG����Q�	���B��q]���B�p�	�������F��IԽ'PN�혪�c����!�:"�[;��:����W���O�P   P   ;$ƽ�4G��ϼ�Aw,��A��xK̿J'̿���,��c����F���Žj�0�4�u��Ù�Ӑ�;�U�;Z����v�]1�P   P   f���k+�Mା�c,����4���C�����Ҫ�,�����"+���|
����&�;���;�ʃ;������P   P   +LZ�Xm��������	�$&�����Rz��>z�������p�	�d��>7���Z�W�����:	�<��<Ӵ�:�ֆ�P   P   ����*��H%6��Ỿ}�B��%̿�C��Rz���C�I'̿��B��⻾<(6��2������<�8�<Q`R<Ȣ<�;�P   P   �x�-�!bؽd� ���B]��%̿��4�wK̿�q]�H���Id���ؽ��-�����z<��z<��z<Z�<P   P   �Z�;�i��WX�����}v���}�B�$&������A����B����7�v�E}����X��Zj����;*m�<��</��<P   P   	��<H��;\y���h����d��Ỿ��	��c,�Aw,�Q�	�O0����d�����vi�g��q�;�g�<7�<��<P   P   �l�<��<E�;\y���WX� bؽG%6�����Mା�ϼ����������6� ٽ�1Y�����Ϡ�;���<KD�<���<P   P   ���<��<��<L��;�i�w�-��*��Vm���k+��4G��KG�,�+����������L.�!>k��͚;���<a�<���<P   P   �;0<�2<���;�8.#'��ͼ�-8�����M��V`�����ὢ����e��i�8�B�μ7�(�_��Ƽ�;�<P   P   �<�<��<jح;�[8����|��TJ���:�;!k�,փ�3䃽�ok��;�����<���"�$!��D��;m�<P   P   ɼ�;W��;&�;w��;�J;��,���ʻ�Z�X6�����l�.R��=���H���|[�y�̻/�8�%�H;E��;P   P   �[��ZR��$J��=�5W �7T.��+#�b6������Eg�����z���~Ȥ��ܒ���g�b��Ţ����%�*�8�^��P   P   5�(���G�5�S��dG��'�NK�G˻:*��Iλ�����$���?�hqJ�i�?���$�K��DϻƢ��y�̻�"�P   P   B�μ����k�����}y���Eμ[���S�Y�2������S��S0������z\�����K�c��|[��<��P   P   i�8�DBp�Gy�������P��(�o��68��2�)��f��J$���e���@���B��{\���$���g�I������P   P   �e����½*���_�
�%�
������}½0�Y:�y��E���S?��|�����@�����j�?��ܒ��켿;�P   P   ����"7���A�h�m���~��Hm��DA���� ��"�j�Y���+����I��|�e����iqJ�Ȥ��=��ok�P   P   �5�6�\��{���\;�s�j������VT6���ws��`���+���S?���S0���?�{���/R�4䃽P   P   ��#Q�P��V��/n<��BU��1<��M��⭾@�P�R��ws��Y���E���J$��S���$�����m�-փ�P   P   W`��Q�]8���'�$���ڿ�����U��U9'��˼�?�P���"�j�y뼀�f��������Eg����<!k�P   P   �M��ˠ6��-���'����=r���3�F�=֡�U9'��⭾VT6� ��Y:�*�3��Kλ���Z6����:�P   P   ���~�������o�_{��Bj���d��d�F��U���M��������0󋽉2�U�Y�<*��e6���Z�UJ�P   P   �-8�<{½�GA��o���9<�ɿ����3���d���3�����1<�j���DA��}½�68�\���K˻�+#���ʻ�|��P   P   �ͼ|o�fT���m���߾�U�ɿ��Bj�<r�ڿ��BU�s྇Hm�����(�o��EμQK�(T.�ɶ,����P   P   /#'��������p
���~���߾�9<�_{�����#���/n<�[;���~�%�
��P��y���'�(�7ܽJ;�Y8P   P   ��8PF�DV�&��p
��m��o���o��'��'�V��z���g�m�_�
���������dG�Z��5r��;gح;P   P   ���;"o�rNR�CV����fT���GA������-��]8��P��[����A�)���Gy��k��7�S�P%J�"�;��<P   P   �2<�v�;o�PF�����|o�;{½~��ˠ6��Q�#Q�5�6�"7���½DBp�������G��R�S��;�<P   P   ����-̻�D���`xӼ�$�!3p��v����н��2���zD�g�н�Ȥ�O�p���$��1Լ9���A���̻P   P   �̻�m̻����5.����T���,�	��;��o�b��-��;���D���p�o�;���	�F<��ř��Q�.�?���P   P   @��������C].��pP��Ʉ�$z��m����x+�˩?��G���?��+�����e�c���A���*Q�Q�.�P   P   8���Y0�����gR��GB���Մ�hZ��D���n��� �߼w���������2���߼^i��np��ѐ��A��ř��P   P   �1Լ��1
꼩��C�Ӽ���������aɤ��N��<k��"����ļ���W���ˢ��3��np��b��E<��P   P   ��$��<�O
J�3�I�0�;��7$���	��������8��SN��Cp��<�� ���董�ˢ��^i���e伤�	�P   P   O�p�	В�3Ѧ�(J��g��������2p�hq;��n��L߼�<��&[��9���7��������V����߼���o�;�P   P   �Ȥ��~׽���[,������F׽X��'Zo��-+��������롼�甼7���������2���+��p�P   P   g�нi'�J�A� �g�ew���g�gA����;н�׍�=?�-V��Aļ�롼9���<���ļ�����?��D��P   P   zD��8�R���6��$̾<̾ծ��A��ؓ7���$˚���F�-V����%[��Bp��!������G�;��P   P   3���!O����d���# �
c2�|��B-񾷽��j�N��-��$˚�=?�����<��RN��;k��v���˩?�-��P   P   ��O���������b�Mϓ�B����Nb���� ��i�N���׍��-+��L߼�8���N���߼x+�b��P   P   ��н��7�~�����瀿��˿�0��)�˿���������ؓ7��;н'Zo��n����`ɤ�m������o�P   P   �v�����a��.m�5�b�L�˿���J��(�˿�Nb�A-�A����X��iq;������D���m���;�P   P   !3p�T׽(pA�_ா ��Ó�,?������0��B���{��ծ�gA�F׽�2p���	����hZ��$z��,�	�P   P   �$��s����a�g��˾rP2��Ó�L�˿��˿Mϓ�
c2�<̾�g���������7$������Մ��Ʉ�T���P   P   `xӼ�;�)q��.����v��˾ �5�b��瀿��b��# �$̾ew���g���1�;�C�ӼHB���pP����P   P   ���R��I�-���.��a�g�_ா-m�����d��6�� �g�[,�(J��4�I����hR��D].��5.�P   P   �D�_����`��I�)q����'pA��a��~���������R���I�A����3Ѧ�O
J�2
����������P   P   -̻�x�_����R��;��s��T׽����7�
O� O��8�i'��~׽	В��<���Z0������m̻P   P   �9��������Ǽ6���ix"�w�W�i��������ڽx��w����f4۽�A���L��SX�-�"�[S����Ǽ¬�P   P   ¬������ʷ���ϼ7������u�>�-�k�V����x��3ի��᫽����� ���'l�JR?�K4�M��Jм,��P   P   ��Ǽ�Mż3�Ǽ��ϼ��l�� 	���'�,B���Z�o)l���r��Kl��Z��SB��(��T�������JмP   P   ZS�������������u���Uw�����:
����ft"�bf-���3���3���-�Ш"���~
�������M��P   P   -�"��L*��-�b.*���"�4��h	��5
�+T���	��1��R����Ze�9V�3
����~
��T�K4�P   P   SX���m���z���z� �m���W���>�i�'����%�	��H�v� �@\���m��� ��s�3
����(�IR?�P   P   �L���O�������f�����Q��Ĝk��A��P"����v �HO�����8q��� �9V�Ш"��SB��'l�P   P   �A��uc��o��R�7C�1G�>��ٴ��Ȍ��8Z�D,-��*�a.���𼰧�m��Ze���-��Z�� ��P   P   f4۽9���8�c�V��gb�nV���7�����ڽ�4��m�k��~3� b�`.��GO��?\�������3��Kl�����P   P   ����,0��}p�q������愭�(>���p���/�5���x��c'r��~3��*��v �u� ��R���3���r��᫽P   P   w�r�B������Ⱦ|)��o$	�����!�Ǿ�>���MB�!� ��x��m�k�C,-����H��1�af-�n)l�3ի�P   P   x��/�B�CĘ�y��9�$��ML��2L���$��d�lx���MB�5���4���8Z��P"�$�	���	�et"���Z��x��P   P   ��ڽ�0�1w����辘�6��#���s�����j�6��d��>����/���ڽ�Ȍ��A����+T����+B�U���P   P   ����R���Ap�L�Ǿ>�$�:"��z���iz�������$�!�Ǿ�p���ٴ�Ük�i�'��5
�:
���'�-�k�P   P   i������7��K��"��kFL��|��z����s���2L�����(>����7�>��Q����>�h	���� 	�t�>�P   P   v�W�W����:�]V��y��r	�kFL�:"���#���ML�o$	�儭�nV�1G������W�4��Tw���l�����P   P   ix"��m��:��"�$8b��y��"��>�$���6�9�$�|)�������gb�7C��f�� �m���"�u����7���P   P   6�����)�:3z��Ƚ�"�]V��K��K�Ǿ���y�辖Ⱦq��c�V��R������z�b.*������ϼ��ϼP   P   ��Ǽ�S��a�,�;3z��:���:���7��Ap�1w��CĘ������}p��8��o�O�����z��-�����3�Ǽ�ʷ�P   P   ����iż�S����)��m�W�����R���0�/�B�r�B��,0�9��uc����m��L*������Mż����P   P   f��Q��}���i0���R��܀���������ݽx���)��B�����ݽ㾽�Q�� ���S���0������P   P   �����YK�l��r0��J�	�k����������� e��(p��B���ќ�+H��6�k��fJ�N0����h�P   P   ����{�������;%��%1���A�odV���l��Ā�Z1���슽�@������m�p�V�pB�;j1�rs%���P   P   ��0�6<1��/1���0��0��)1���4���;��E��`O��AX�<u]���]�7eX���O��^E��<�U05�;j1�N0�P   P   �S���Y��0\���Y���R�J���A���;�p�8�W�8�3�:��~<�*O=���<���:�b9�"9��<�pB��fJ�P   P   ��၊��󏽲菽�b��H䀽g�k�~TV�E�2�8��`1��}-���+�D�+�.�-�7�1�b9��^E�p�V�6�k�P   P   �Q���X������aƽ�����!��F��\��'�l��<O� �:��p-�Qt&�6N$�!�&�-�-���:���O�m�*H��P   P   㾽g0㽲i���
�,�
�H����݆�����v����X��V<���+��C$�5N$�D�+���<�7eX������ќ�P   P   ��ݽ=��zd)�C&@��H��@�e))����
uݽ����l����)]�n=���+�Pt&���+�)O=���]��@��A��P   P   B����W#�2S�k4��3����w����)�R��#��:��������)]��V<��p-��}-��~<�;u]��슽(p��P   P   )���^1��t�㟾5C��'Z;���6���I�s��1�-�����l����X��:��`1�2�:��AX�Z1���d��P   P   x���T1�ds��F�����쾠�	���	��c��?��<���1��:������v����<O�2�8�W�8��`O��Ā�����P   P   �ݽ'<#�ot�w|���"����#���3���#�?����?��I�s��#�
uݽ���'�l�E�o�8��E���l����P   P   ��������R�nϟ�ܖ�H�#��eG��XG���#��c�6���)�R����݆��\��~TV���;���;�ndV����P   P   �����⽱7)�����0��U�	���3��eG���3���	������e))����F��f�k���A���4���A��k�P   P   �܀�T��zA�c�?��s��wV;U�	�H�#���#���	�'Z;�w���@�H��!��H䀽J��)1��%1��J�P   P   ��R��L��%���N�
�ߩH��s���0��ܖ쾳"�����5C��3����H�,�
������b����R��0��;%�q0�P   P   �i0��rY��Ï��,ƽN�
�c�?����nϟ�w|��F���㟾k4��C&@���
��aƽ�菽��Y���0����l��P   P   }���1�m�[��Ï�%���zA��7)��R�ot�ds���t�2S�zd)��i�����󏽟0\��/1���XK�P   P   Q���\��1��rY��L��T��������'<#�T1��^1��W#�>��h0㽐X��၊���Y�6<1��{����P   P   
o8�"D<�>H�L\���z��;���^��C�ý�۽T������Bܽ9�ýϏ���g����z���\�#+H��V<�P   P   �V<�M<��QA�	�K��H\��s��ˇ�痽|᧽�������(������a��������PXs�T�\���K��nA�P   P   #+H��F�"H���K��R��N]�@�k�=}��܇��^��Ek��\����x���w��h����_}���k��]�e�R���K�P   P   ��\�� ]��]�k�\�tR\��P]�*k`���e��nm���u��|��a���g��p�|���u�?�m��:f��`��]�T�\�P   P   ��z��;���A���-���z��s���k�T�e�/�b���a�Fcb��kc�;�c���c��b�� b�_�b��:f���k�OXs�P   P   �g��HF��cŝ�p����*���?���Ǉ�#}��]m��a�
Z���U�*�S���S�b�U�pFZ�� b�>�m��_}����P   P   Ώ��ҹ�&�Ž��ɽvgŽ����V��֗��ɇ��wu�"Kb�£U���N��[L��N�b�U��b���u�g������P   P   9�ý�Q�S����Y��O�;d��R	ཞkýؾ��>��]s|�	Ec�ıS��PL��[L���S���c�o�|��w��`��P   P   Bܽ�?�����2*�QB0��*�/�����۽�̴�|=���>��t�c�ıS���N�)�S�:�c��g���x�����P   P   ��A��9q7��%V�y�h�Y�h���U��07��G�_9��:���i���>��Ec�£U���U��kc��a��\���'���P   P   �����+�M�4�~��$���˚������~���M�ui�̩��:��|=��]s|�!Kb�	Z�Ecb��|�Ek������P   P   S������V�=&���w��=s��Yd���R������_6V�ui�_9��̴�>���wu��a���a���u��^�����P   P   �۽�r�!�M��!��>����۾�����ھ_Y��������M��G��۽ؾ���ɇ��]m�.�b��nm��܇�{᧽P   P   C�ý%�%V7���~��q��N۾ش��ܨ����ھ�R����~��07����ký֗�"}�S�e���e�<}�痽P   P   �^��z�����V�t��&t����ش�����Yd�������U�/��Q	ཐV���Ǉ���k�)k`�@�k��ˇ�P   P   �;��睹��^��*���h� ̚�&t��N۾�۾=s���˚�Y�h��*�;d������?���s��P]��N]��s�P   P   ��z�����PŽA�800���h�t���q��>����w���$��y�h�QB0��O�vgŽ�*���z�tR\��R��H\�P   P   L\����힝�U�ɽA�*��V���~��!��=&��4�~��%V��2*��Y���ɽp����-��k�\���K�	�K�P   P   >H���\�"&��힝��PŽ�^�����&V7�!�M���V�+�M�:q7����S���&�Ždŝ��A���]�"H��QA�P   P   "D<���F���\�������睹�z�%��r�������B���?��Q�ҹ�HF���;��� ]��F�M<�P   P   Ta��ud�5�n��j���4��d������Y�Ž8!ؽ<U��(�_e� ?ؽo�ŽC��9ܝ�oT��@����o���d�P   P   ��d�,~d�%i��[r�:`��z�������+��������ȿ�sп����ׯ�\)��G���6��|�� �r�� i�P   P   �o�|�m���n��br��}x�)Հ��ꆽC"��t���Q����S��+���_��I����Օ�mC��D���󀽜�x� �r�P   P   @���墀�w����s���c��|Հ�W���W���P��j����G��'⎽R玽�W��h���jn���x��W=����|��P   P   oT��O���"u��2���<��+���膽@U��s���������<��O`��+F������$ӂ��x��D���6��P   P   9ܝ�	6��ͧ��ħ�z��P���k약���TH�������|�hRx��Vv��`v�px�D�|���jn��lC��F��P   P   C������ǽ�\ʽǽ�齽�������˦��]v����aFx�g�q�|}o�c�q�px���h����Օ�\)��P   P   n�Ž-�۽���(��Q���s���X۽'sŽ֛��Wl���/���)��I?v�Vro�|}o��`v�+F���W��H����ׯ�P   P   �>ؽ�X��TA��������l �7��U�׽dй�*,���8H��I?v�g�q��Vv�O`��Q玽�_����P   P   ^e彇	�Ե ��+5��BA�6A��	5�{� ����9��ᢽ��)��`Fx�hRx�<��'⎽*��rп�P   P   �(��F���/�V<O��>g��Op�n!g��O��/���N���*,���/���󁽽�|�����G���S���ȿ�P   P   ;U影A��l5�}�^�x_��������lI���^��75���9�dй�Vl��]v��������i���P�������P   P   8!ؽ�	���/���^�&��ԣ��z@��}���쇾�^��/����U�׽֛��˦��TH��r����P��t���*���P   P   X�Ž3��c� �e/O��\������w������}���lI���O�{� �7��&sŽ�������@U���W��C"�����P   P   ���<h۽E,��5��5g�����F��w���z@������n!g��	5�l ��X۽���k약�膽W���ꆽ��P   P   d����载"����R8A��Rp��������ԣ�����Op�6A���s���齽O���+��|Հ�)Հ�y��P   P   �4��@����ƽ������S8A��5g��\��&��x_���>g��BA����Q���ǽz��<���c���}x�:`��P   P   �j��H���G����Aʽ�������5�e/O���^�}�^�V<O��+5���(���\ʽ�ħ�2����s���br��[r�P   P   5�n�ǎ�� _��G�����ƽ"��F,�c� ���/��l5���/�Ե �TA�����ǽͧ�"u��w�����n�%i�P   P   �ud���m�ǎ��H���@���载=h۽3���	��A��F��	��X��-�۽���	6��O���墀�|�m�,~d�P   P   Nv�����r��`�����|	��+R��jƽ�ӽ��ݽ+/�ηݽ]Խ�ƽq���'��Ǚ�c��������P   P   ���U���G�򈽤���%���͠�%7��K ��B��
j���o��!���8��T��u렽�B��6&�����+���P   P   �������gx��P���z���ey��5���ie��ht���ҥ�����窽D���x好L���c�������Д���������P   P   b��;-��{(��J�����ay������`M�����<"��U@���|��J���_N���7��ٻ��`k��v���Д��6&��P   P   Ǚ�o���A��ύ�������&��j����J��ɐ����^ҏ����<�4鏽�㏽����搽`k�������B��P   P   �'���+�����������	���Ǡ��]�����=���������뽉�������>ь����ػ��c���u렽P   P   q���P���0ǽ�ɽ'ǽ'1���H���(��9d��=���Ǐ�����'������h��������㏽�7��K���T��P   P   �ƽq�ֽ��㽍Y�KN�8�㽌dֽ��Žz�������*���Ϗ�>���x��������4鏽^N��x好�8��P   P   ]Խ2P�C:��	�j��	�B"�,��ӽ�޼�4k��j`��}ۏ�>���&���꽉�;�I���C��� ��P   P   ͷݽ���O����h�$���$�K�� /������wݽ�:�����j`���Ϗ�������������|���窽�o��P   P   */���=l���-�բ<��#B�@�<���-�G�&������:��4k���*���Ǐ����]ҏ�T@�����	j��P   P   ��ݽ����z7��RN�M�[���[��7N��V7�>��&���wݽ�޼�����=��<�����;"���ҥ�B��P   P   �ӽ�����e�Cx7���T��#k��{s��k�#�T��V7�G������ӽz��9d�����ɐ����gt��J ��P   P   iƽ5��C��-��PN�%k��q|��j|��k��7N���-� /�,���Ž�(���]���J��_M��he��%7��P   P   +R���rֽ2,�����<�#�[��s��q|��{s���[�@�<�K��B"��dֽ�H���Ǡ�j�������4����͠�P   P   {	��g2�����h	���$�K'B�#�[�%k��#k�M�[��#B���$�	�8��&1���	���&��`y��ey���%��P   P   �������ǽ�C뽕����$���<��PN���T��RN�բ<�h�$�j��KN�'ǽ���������z������P   P   `��o���8ᮽ��ɽ�C�h	����-�Dx7��z7���-�����	��Y��ɽ��ύ��J��O�����P   P   �r�����0��9ᮽ�ǽ���2,��C��e��>l�	O�C:���㽭0ǽ����A��{(��gx��FP   P   �񂽭������o������h2���rֽ5������������3P�r�ֽ�P���+��o���;-������U���P   P    ^������_��c����D��z孽�Ĺ���ŽP	н�)׽\�ٽO3׽�н
�Ž�ܹ�����Z��޳��l��Y���P   P   Y��������J������൚��F������~&��ʸ�nǾ�*½�½�Ӿ��ݸ�:>�����_���ʚ�Թ���T��P   P   l������Dd��g���-嗽]���-��ۣ�R���ɬ��������h����ج������ G��/��G���Թ��P   P   ޳������L���i���x���!����Y���&�����(���`�������>���� ��#>��Hs�����/���ʚ�P   P   
Z��~Ĥ��E�������G���F���*���V��{��9J��b�����������������`��{"��Hs�� G��_��P   P   �����ᱽ#��#���б�T䭽����2ԣ�a���F���q��쥖�8̕�}Е�Ҳ�������`��#>�������P   P   �ܹ�^_��C�ƽJ[Ƚozƽ�E��������!����������c�������<��a��Ҳ������ �����9>��P   P   	�Ž&�ѽX�۽����,�۽,�ѽ��Ž|�����������X㚽���7���<��}Е�����>����ج��ݸ�P   P   �н��ὥ��xy��72 ��e��mb�$�὘�Ͻ𨾽y���D~���ᚽ�����8̕���������h����Ӿ�P   P   O3׽�d��}���2��X��٘�g�2��׽�������D~��X㚽b���륖���`��������½P   P   [�ٽ�g��DP	�r��� ���#�u �ȋ�66	��3��҈ٽ���y������������q��b���'������)½P   P   �)׽�c�����.��e+��93�33�. +�J��ǫ��3���׽𨾽��������F��9J�����ɬ�mǾ�P   P   O	н�W�L	����/��E<��A��:<���.�J��66	�2�Ͻ|��� ���a��{���&��R���ʸ�P   P   ��Ž?�Ὁv�����+��F<�@F��;F��:<�. +�ȋ�g�$�ί�Ž���1ԣ��V��Y��ۣ�}&��P   P   �Ĺ���ѽ�r񽣢�� ��;3�h"A�@F��A�33�u �٘�mb�,�ѽ��������*���󛽪-������P   P   y孽nH����۽�j��|��]�#��;3��F<��E<��93���#�X���e��,�۽�E��T䭽�F��!��]���F��P   P   �D��e̱��tƽ�
�O/ �|��� ��+�/�e+�� �2��72 ���ozƽ�б��G��x���-嗽ߵ��P   P   c���1������&NȽ�
��j�����������.��r����yy����J[Ƚ$������i���g�������P   P   �_�������8������tƽ��۽�r�v�L	����DP	��}����X�۽C�ƽ#���E��L���Dd���J��P   P   �����������1���e̱�nH����ѽ@���Wc���g���d����&�ѽ__���ᱽ~Ĥ�������������P   P   ̟������򵞽:ģ������첽���S�Ľy�̽�ѽl�ӽ&�ѽ��̽�
Žs�� ��2����ң�������P   P   ����������ʟ��ޣ�B��!$���p���B��ÿ��=½[A½Ϳ� R������8��	.��w�؟����P   P   �����a�������˟�,����7���v��a��pή������+��8���K2���
���߮��3��D����K��<���؟�P   P   �ң�*̣�Wȣ��ǣ��ߣ�%7��w뤽 ���`��fΨ����E���������/ި�u���������K��w�P   P   2���{ë�$��U���Ρ��J��Tt��s����礽�;���磽Ṭ�1ɣ�kӣ�g����N��8������D���	.��P   P    �����畷����3赽벽������Z��[8���ޡ��V���������{a��𡽴N��u���3��8��P   P   s������l�Žh�ƽt�Žf��������e���®��è��ߣ�fR���/���{��h7��{a��f���.ި��߮�����P   P   �
Ž1νV-սtٽ�ٽ�ս��ͽ��Ľ�0��챽��E���l����w���{�����kӣ�����
�� R��P   P   ��̽��ٽ����o�(�Xa�P�佞vٽ��̽�������H���i���l����/������0ɣ����K2��Ϳ�P   P   &�ѽ#��&Z����$��*��;���T9�*m��ѽ}½|ش�H���E���fR���V��Ṣ�E���7���ZA½P   P   k�ӽ3������h�����"����b��Ј���_�d�ӽ}½����򩽛ߣ��ޡ��磽����+���=½P   P   �ѽE��%����
�����	��q��B�
�����_��ѽ����챽�è�Z8���;��fΨ�����ÿ�P   P   x�̽��p�����
�yr���ے!�����e�B�
�Ј��*m⽣�̽�0���®��Z���礽�`��oή��B��P   P   S�Ľ<�ٽ�P򽱺����g���$�>�$����q��b��T9�vٽ��Ľ�e����s���~ ��a���p��P   P   ����νպ�&���F������!��$�ے!�����;���P����ͽ�������St��w뤽�v�� $��P   P   �첽r���սuf����g%���g�����	��"�*��Xa��սf���벽J��%7���7��B��P   P   �����嵽k�Ž�ٽ�%����F�����yr������$��(��ٽt�Ž3赽Ρ���ߣ�,����ޣ�P   P   :ģ�X���0�����ƽ�ٽuf�'��������
���
�h������o�tٽh�ƽ���U����ǣ��˟��ʟ�P   P   򵞽<���4��0���k�Žսպ佌P�q���%������&Z���W-սl�Ž畷�$��Wȣ��������P   P   ����[��<���Y����嵽r����ν<�ٽ���E��3��#�⽊�ٽ1ν�������{ë�*̣��a������P   P   ɞ��Gq���妽檽pC�����������<Ľ��ɽӴͽ�Ͻ�ͽ/�ɽIĽP���y���sQ���񪽀��u��P   P   �u��s��А��yǧ����|���ǳ���������[T���*½�-½4\��� �������׳��/������ҧ�3���P   P   ��`���I覽hȧ�xC��CS���ܭ������~���浽Ȋ�����e���t����\�����c���Q���ҧ�P   P   ��G窽�㪽�誽E���R���૽s���í��Ԯ�ܶ��w8���;������ᮽ�ӭ� ˬ����c�����P   P   sQ��c���c�����D��+���ڭ������ԫ��A���񪽱Ϫ�H˪��ժ������Q���竽 ˬ���/��P   P   y����︽�%���!��\丽����,ó�����4����>��mW�� ���t��qw��,���e���Q���ӭ�\����׳�P   P   P�������|�Ľ��Ž��Ľ����ރ��y���u���ˮ�z몽|���S���¥��Z��+�������ᮽ�������P   P   IĽ��ʽ�н��ҽ�ҽ�н��ʽI0Ľ5漽9ص�ȩ���Ū��m��z����¥�qw���ժ����t�� ��P   P   /�ɽ�Mӽ�G۽Ȭང�⽾��/4۽4ӽ�ɽ�@���w���'��d����m���S���t��G˪��;��d���4\��P   P   �ͽ �ٽ*�佫s�-�-(�cc�߻�t�ٽͽ�½X���'���Ū�|�� ���Ϫ�w8������-½P   P   �Ͻ>ݽ�L�cg��P����K�f���+R���1�=!ݽ��ν�½�w��ȩ��z몽mW����ܶ��Ȋ���*½P   P   Ҵͽ�;ݽy�����'r������Uj�p����|�=!ݽͽ�@��9ص��ˮ��>���A���Ԯ��浽[T��P   P   ��ɽY�ٽI�_������W�7��R���p����1�t�ٽ�ɽ5漽u��4����ԫ�í��~������P   P   �<Ľ�Cӽ����c��r�>X��+��)��R�Uj�+R��߻�4ӽI0Ľy�����������s�����������P   P   ������ʽ�>۽�n�˫��v���9��+�7���f���cc�/4۽��ʽރ��+ó��ڭ��૽�ܭ��ǳ�P   P   ���������н����,�N�v��?X��W�����K�-(򽾡��н��������+���R��BS��|��P   P   pC��㸽H�Ľu�ҽ]���,�˫��r���'r�P����-򽄒��ҽ��Ľ\丽D��E��xC�����P   P   檽���,����Žu�ҽ����n��c��_�������cg���s�Ȭ���ҽ��Ž�!������誽hȧ�yǧ�P   P   �妽�ު�D\��,��H�Ľ�н�>۽���I�z��L�*���G۽�н}�Ľ�%���c���㪽I覽А��P   P   Gq��񚦽�ު����㸽������ʽ�CӽZ�ٽ�;ݽ>ݽ �ٽ�Mӽ��ʽ�����︽c��G窽`���s��P   P   ����f��S���q�����s��蠾���ý<�ǽ#�ʽ��˽Ǌʽ��ǽӡý���n~��b����z��Y��i��P   P   i���g��J���	��ڐ��G����I���麽0������c½�½����79������W��4ǳ��������O��P   P   Y�����U��@
���7���Ұ�zȲ��𴽣���ݸ�������T���渽���m����ֲ�Bఽ�C�����P   P   �z��Dn���k���s��%���8Ұ�:D��鱽�����z�����z~�������&������[���`����S��Bఽ���P   P   b����5��Vi���0������츳��Ʋ��籽�5��ջ���t���R��K���W���~���Ȱ��E��`����ֲ�4ǳ�P   P   n~���&��-���������p��F��촽ͪ��&����4���1������E���I9��-A���Ȱ�[���m���W��P   P   ���X���I�ý�ĽN�ý�������h⺽���s���o���.��xͬ��W��GӬ�I9���~�������������P   P   ҡý�Ƚg<̽�?ν?<ν�1̽�sȽ�ýM$��xҸ�&��KJ��۪��U���W��E����W���&���渽79��P   P   ��ǽ�νdLԽ�ؽ�rٽKؽ�=Խ��ν��ǽ�������p��@��۪��xͬ�����K������T������P   P   Ǌʽ#5ӽ�۽��zW�oS��ὧ�ڽ�ӽ�tʽ����t���p��KJ���.���1���R��z~������½P   P   ��˽�ս{�߽��������Z���罩�߽�սgl˽�������&���o���4���t��������c½P   P   #�ʽ�ս�.�A����3��2/����󽝠���ս�tʽ���wҸ�s��&���ջ���z���ݸ�����P   P   <�ǽN0ӽ�߽������������e��"���������뽩�߽�ӽ��ǽM$�����ͪ���5���������0��P   P   ��ý�ν#۽����������� ��� �"�������罧�ڽ��ν�ýh⺽촽�籽鱽���麽P   P   蠾�-{Ƚ�EԽ��֑��5�� i��� ��e��2/��Z���ὒ=Խ�sȽ���F���Ʋ�:D��zȲ��I��P   P   s��,���C5̽�ؽ�W����5����������3�����oS�Kؽ�1̽�����p��츳�8Ұ��Ұ�G���P   P   ���*����ý�;ν-rٽ�W�ב������������zW��rٽ?<νN�ý�������%����7��ڐ��P   P   �q���-��4��ؔĽ�;ν�ؽ�ὤ�罘��A�뽶���ὦؽ�?ν�Ľ����0���s��@
���	��P   P   S���g���c��4����ýC5̽�EԽ#۽�߽�.�|�߽�۽dLԽh<̽I�ý-��Vi���k��U��J��P   P   f������g���-��*��,���-{Ƚ�νO0ӽ�ս�ս#5ӽ�ν�ȽX����&���5��Dn������g��P   P   �V���װ�SV��A����㷽f���cm���ý%ƽ�*Ƚ��Ƚn-Ƚ�*ƽo!ý�u��B����췽�Ĵ��[���ڰ�P   P   �ڰ��ذ����u岽Hش�1B��P�'����������/������L���� ��t��� ���zL��[ᴽ�첽����P   P   �[��)��X���岽�ϳ��������*/���Ź�������OX�����p$��)Ϲ�:���������qٳ��첽P   P   �Ĵ�Ҷ��紴�����cش����h��p㵽�v����������˷�_ͷ��������䁶��ﵽ�t�����[ᴽP   P   �췽�Y������ZU��"䷽�@��ˌ��!⵽4Y������J���뜴�����'���´�>��Pf���ﵽ����zL��P   P   B���QѼ�\{���x��Mʼ�\���OﹽM+���s��V���~Ƴ��������;��� ���г�>��䁶�:�� ���P   P   �u��A���bIý��ýDý���~h��(���������:�������)㱽凱��籽 ��´����)Ϲ�t���P   P   n!ý��ƽZgɽ=�ʽc�ʽ_ɽݧƽ�ý������s}�����A���Å��凱�;���'�������p$��� ��P   P   �*ƽ�˽�6Ͻ��ѽ]�ҽk�ѽ�+Ͻ�˽�ƽ�����������ϊ��A���)㱽�������_ͷ����L���P   P   n-Ƚ�nνt	ԽEؽW�ڽ@�ڽ$<ؽ��ӽ�^νMȽi��� J�����������������뜴��˷�OX�����P   P   ��ȽQ:н<׽�ݽ��� S⽰���	ݽA-׽�)нq�Ƚi�������s}��:���~Ƴ�J����������/���P   P   �*Ƚ9нEZؽ��߽�;��<�:�g3�r�߽�Kؽ�)нMȽ���������V�����������������P   P   %ƽ`kν':׽F�߽��潛q����l뽾��r�߽A-׽�^ν�ƽ�������s��4Y���v���Ź����P   P   �ý�˽�Խ�ݽ�;彆r������l�g3��	ݽ��ӽ�˽�ý(���M+��!⵽o㵽*/��'���P   P   cm���ƽ�1ϽCؽ����>�������:轰��%<ؽ�+Ͻݧƽ~h��Oﹽʌ��h������P�P   P   f���w���%bɽ�ѽ��ڽ�U��>轆r뽛q��<� S�@�ڽk�ѽ_ɽ���\����@��������1B��P   P   �㷽�ɼ�Dýo�ʽ�ҽ��ڽ��཭;彋���;����W�ڽ]�ҽc�ʽDýMʼ�"䷽cش��ϳ�Hش�P   P   A���kS��Pv����ýo�ʽ�ѽCؽ�ݽF�߽��߽�ݽEؽ��ѽ>�ʽ��ý�x��ZU�������岽u岽P   P   SV��α���{��Pv��Dý%bɽ�1Ͻ�Խ':׽EZؽ<׽t	Խ�6ϽZgɽbIý\{������紴�X�����P   P   �װ��%��α��lS���ɼ�w����ƽ�˽`kν9нQ:н�nν�˽��ƽA���QѼ��Y��Ҷ��)���ذ�P   P   '�����p5��~���j���*���
��;�½��ĽDqƽ+�ƽ�sƽ��Ľ4�½����1��Cq�����9��9��P   P   9�������������� ���������������ʿ��&�����������*���п���8������[(��U���k���P   P   �9������6�������Y���L���n�����[ֻ�Լ�h~���������Zټ��ݻ�ݱ��/x���U��a��U���P   P   ��J��� ��e	��� ��\L��������]��(ɹ��!��S���T���&��Pй��f�����������U��[(��P   P   Cq��p���uݺ������j���󹽃m����냸��6��I��췽巽X﷽���n?��z�������/x������P   P   �1�����������������(��_�������[��5���M�������]���_������V��n?���f��ݱ��8��P   P   ��������½�?ý�½۸��������1ѻ��Ĺ��������:ֵ�Ґ���ٵ��������Pй��ݻ���P   P   4�½	aŽSVǽ�aȽ|_Ƚ�Oǽ:WŽ˸½�ÿ��̼� ���淽�Y������Ґ���_��X﷽�&��Zټ��п�P   P   ��Ľ��Ƚ��˽�{ͽ�(ν�wͽ߁˽P�Ƚ��ĽE���t��oJ���ݷ��Y��:ֵ��]��巽�T������*��P   P   �sƽl�ʽ6�ν� ҽ��ӽx�ӽ��ѽ��ν��ʽ4fƽ����}���oJ���淽��������췽S����������P   P   +�ƽJC̽�Dѽbdս�ؽ�ٽ�ؽX\ս�9ѽ�6̽��ƽ�����t�� ������M��I���!��h~������P   P   DqƽrB̽�ҽ�6׽�۽�*ݽ�(ݽ�۽�-׽ҽ�6̽4fƽE���̼��Ĺ�5���6��'ɹ�Լ��&��P   P   ��Ľ��ʽlCѽ�6׽o ܽ�`߽`��}]߽9ܽ�-׽�9ѽ��ʽ��Ľ�ÿ�1ѻ�[��냸��]��[ֻ��ʿ�P   P   ;�½��Ƚ��ν�cս�۽�a߽������}]߽�۽X\ս��νP�Ƚʸ½������������������P   P   �
���[ŽD�˽C�ѽ�ؽ8,ݽ��བ��`�འ(ݽ�ؽ��ѽ߁˽:WŽ��_����m�������n������P   P   �*�����kRǽ�yͽ?�ӽٽ8,ݽ�a߽�`߽�*ݽ�ٽy�ӽ�wͽ�Oǽ۸���(����\L���L������P   P   �j�����.�½�_Ƚ<)ν?�ӽ�ؽ�۽o ܽ�۽�ؽ��ӽ�(ν|_Ƚ�½����j��� ���Y��� ��P   P   ~��Z���琾�A=ý�_Ƚ�yͽC�ѽ�cս�6׽�6׽bdս� ҽ�{ͽ�aȽ�?ý��������d	����������P   P   p5�������ٺ�琾�.�½kRǽD�˽��νlCѽ�ҽ�Dѽ6�ν��˽TVǽ�½����uݺ�� ���6������P   P   ��������Z����������[Ž��Ƚ��ʽrB̽JC̽l�ʽ��Ƚ	aŽ�������p���J��������P   P   ����N���,������V���c��K����½Y!Ľ�2Žu�Ž�4ŽT$Ľ��½�����i���[��\���0��\P��P   P   \P��<O��x���2��� ���� ��2���q��V���S�����������V���Z��/	������.��Q���膹�)���P   P   0������-��a�������ĺ�����G���eg��m"��ў���ʾ�����&��Sm��[���t����˺�g��膹�P   P   \���������������2����ĺ�F���A�������޻�p���A��	C��&!��_份���I��h���˺�Q���P   P   �[��E���	���"����V����������>@��#<��������s��Fo��av��򎺽L���{���I��t���.��P   P   �i��.��%l���j�����mb�� ����������������)���BG���H��f���:��L������[�������P   P   ����������½��½w�½ӿ��Y���u����c��ۻ�󆺽�����ḽ����s丽f���򎺽_份Sm��/	��P   P   ��½�nĽS�Ž��ƽ�ƽ1�ŽgĽ�|½�P��J��N���o��VD����������H��av��&!���&���Z��P   P   T$Ľ �ƽ��Ƚ�Jʽ��ʽ�Gʽ3�Ƚ=�ƽ?Ľ0L��~����:���i��VD���ḽBG��Fo��	C������V��P   P   �4ŽkȽb˽�ͽ&�ν�ν��ͽnZ˽�uȽ:*Ž���������:���o������)����s���A���ʾ�����P   P   u�Ž�kɽ�ͽ	�ϽL�ѽ�ҽ8�ѽ�Ͻ�̽:bɽ��Ž����~���N��󆺽��������p��О������P   P   �2Ž%kɽ��ͽ�<ѽ��ӽflս�jս��ӽ�5ѽ�ͽ:bɽ:*Ž0L��J��ۻ����<����޻�m"���S��P   P   Y!Ľs}Ƚͽ%<ѽ�Խ�ֽW�׽e�ֽ��Խ�5ѽ�̽�uȽ?Ľ�P���c������#����eg��V��P   P   �½þƽ`˽��Ͻ��ӽ��ֽ��ؽ��ؽe�ֽ��ӽ�ϽnZ˽=�ƽ�|½u�����>@��A��G���q��P   P   K����jĽ��Ƚ�ͽ��ѽ�mս��׽��ؽW�׽�jս8�ѽ��ͽ3�ȽgĽY��� �������F�������2���P   P   �c������V�ŽzIʽN�ν�ҽ�mս��ֽ�ֽflս�ҽ�ν�Gʽ1�Žӿ��mb�������ĺ��ĺ�� ��P   P   �V�������½�ƽ?�ʽN�ν��ѽ��ӽ�Խ��ӽL�ѽ&�ν��ʽ�ƽw�½����V��2������ ���P   P   ���4����i��P�½�ƽzIʽ�ͽ��Ͻ%<ѽ�<ѽ	�Ͻ�ͽ�Jʽ��ƽ��½�j��"�������a���2���P   P   �,��˄��b����i����½V�Ž��Ƚ`˽ͽ��ͽ�ͽb˽��ȽS�Ž��½%l��	��������-��x���P   P   �N�����˄��4�����������jĽþƽs}Ƚ%kɽ�kɽkȽ �ƽ�nĽ����.��E����������<O��P   P   Z����ź��l���u���˽��Q��1����Y½��ýWOĽ7�Ľ�PĽ�ý�\½c����V��|Ͻ�;y��Io��Ǻ�P   P   Ǻ�(ƺ���]�����������ܭ��mȿ�����wz����������|�������̿�ﲾ������������Z��P   P   Io���W��um��w������֢��(G��+�������n ���z��Ú���|���#��P�������M��w���:�����P   P   ;y��{p��zo��Fv��Ć��|���B˼������:���r��Y�����������8���Gw��J@�����Ѽ�w�������P   P   |Ͻ�������(����˽�ƍ��TF�������¼�����Bs��Qa���[��*c���w��I���Vɼ���M������P   P   �V���п�������Ϳ��P��3���1��8������5
������}��Q��������I���J@������ﲾ�P   P   c��������d½½Ab½L�������9ſ������o��q�������2��	���4�������w��Gw��P����̿�P   P   �\½��ý��Ľ�UŽ0TŽ��Ľs�ýtU½����z��c����]���{�����	��Q��*c��8����#������P   P   �ý�tŽ ǽ�Ƚ,[Ƚ��ǽ��ƽ�mŽ�ý�t��u��.���jW���{���2���}���[�������|���|��P   P   �PĽ?�ƽ��Ƚ.Wʽ�)˽�'˽Sʽ��ȽۮƽIĽz���哿�.����]���������Qa������Ú�����P   P   6�Ľaǽ��ɽI̽�pͽ��ͽ�nͽ�̽�ɽ�Yǽq�Ľz���u��c���q��5
��Bs��Y����z������P   P   WOĽj`ǽ�^ʽx�̽G�ν��Ͻ��Ͻ��νE�̽�Xʽ�YǽIĽ�t��z���o�����������r��n ��vz��P   P   ��ý޴ƽ
�ɽ8�̽osϽ�ѽj�ѽ�ѽpϽE�̽�ɽۮƽ�ý���������8���¼��:����������P   P   �Y½rŽ�Ƚ�̽t�ν'ѽ�/ҽ/ҽ�ѽ��ν�̽��Ƚ�mŽtU½9ſ�1���������+���mȿ�P   P   0���9�ý��ƽsVʽ`qͽ��Ͻ��ѽ�/ҽj�ѽ��Ͻ�nͽSʽ��ƽs�ý����3���TF��B˼�(G��ܭ��P   P   �Q��������Ľ� Ƚ�)˽�ͽ��Ͻ(ѽ�ѽ��Ͻ��ͽ�'˽��ǽ��ĽL����P��ƍ��|���֢������P   P   �˽�NͿ�pb½�TŽ�[Ƚ�)˽`qͽt�νosϽG�ν�pͽ�)˽-[Ƚ0TŽAb½Ϳ��˽�Ć���������P   P   �u��V��������½�TŽ� ȽsVʽ�̽8�̽x�̽I̽.Wʽ�Ƚ�UŽ½���(���Fv��w���]���P   P   �l��n��O�����pb½��Ľ��ƽ�Ƚ
�ɽ�^ʽ��ɽ��Ƚ ǽ��Ľ�d½�����zo��um����P   P   �ź�+V��n��V���NͿ�����9�ýrŽ޴ƽj`ǽaǽ?�ƽ�tŽ��ý�����п�����{p���W��(ƺ�P   P   �u��"������k佽u㾽���y.��A@½qý��ý��ý�ý� ý�B½�1��	��y澽%罽���0���P   P   0���v���ݼ�bP��5󽽪�������O]�����ϛ��&���������������`�������������9S��߼�P   P   ���������\P��頽��	��惾�����|���߿��!��^8��;#��n⿽����;	��|���_������9S��P   P   %罽W߽�T޽��佽>󽽻	��)���O��z����������Ӿ��Ӿ��þ�D����~���T��4.��_�����P   P   y澽���p�����@㾽������CO��6!������㽽tԽ�=Ͻ� ֽ�W潽a ���&���T��|�������P   P   	��Pb������Đ��N_�����`���M���x�����c���[N��*��A+��&Q��h���a ���~��;	������P   P   �1�������G½m½�E½����v,���Z��?z��f���`ώ�M��}�kѼ� �&Q��W潽D��������`��P   P   �B½4Gý�ĽAmĽlĽ�ĽiBý7=½���&ܿ�i����ѽ�C(��Kм�kѼ�A+�� ֽ��þ�n⿽���P   P   � ý˄Ľ�Ž�_ƽt�ƽ^ƽ�Ž�Ľ)ý,���6���ξ��˽�C(��}�*��<Ͻ��Ӿ�;#������P   P   �ý�mŽ��ƽ�Ƚ��Ƚg�Ƚ�Ƚj�ƽ5hŽ�ý����3���ξ��ѽ��M��[N��tԽ�Ӿ�^8������P   P   ��ý#�Ž��ǽ�Nɽ�IʽƠʽ�GʽKɽ��ǽ��Ž��ý����6��i���`ώc���㽽�����!��%���P   P   ��ý��Ž�Ƚ�ɽ�Z˽�̽�̽8X˽Q�ɽ
Ƚ��Ž�ý,���&ܿ�f���������������߿�Λ��P   P   qý�lŽ#�ǽ�ɽ˹˽��̽�CͽA�̽��˽Q�ɽ��ǽ5hŽ)ý���?z���x��6!��z���|�����P   P   A@½�Ľ��ƽ9Nɽ�Z˽��̽o�ͽ��ͽA�̽8X˽Kɽj�ƽ�Ľ7=½�Z��M��CO���O�����O]��P   P   y.���Dý��ŽVȽ�Iʽk̽Eͽo�ͽ�Cͽ�̽�Gʽ�Ƚ�ŽiBýv,��`������)��惾�����P   P   �������ĽJ_ƽ��Ƚ�ʽk̽��̽��̽�̽Ơʽg�Ƚ^ƽ�Ľ�����������	���	������P   P   u㾽�_���E½slĽ�ƽ��Ƚ�Iʽ�Z˽˹˽�Z˽�Iʽ��Ƚt�ƽlĽ�E½N_��@㾽>�頽�5�P   P   k佽 ������Xl½tlĽJ_ƽVȽ9Nɽ�ɽ�ɽ�Nɽ�Ƚ�_ƽAmĽm½Đ������佽\P��bP��P   P   ���aݽ�5�������E½�Ľ��Ž��ƽ#�ǽ�Ƚ��ǽ��ƽ�Ž�Ľ�G½����p��T޽����ݼ�P   P   "���o��aݽ� ���_������Dý�Ľ�lŽ��Ž#�Ž�mŽ̄Ľ4Gý����Pb�����W߽����v���P   P   d佽9��+b������=���r���Fg���0½[�½�<ý�`ý;=ý�½3½�i�����ٷ��)����c����P   P   ��y��b1��ӈ��k�������2������S���������Z���k���0U������%6��͘��-�����3��P   P   �c���V���b��ӈ���ľ�����o���Ϳ�{'��-p�����v������Mr���*��5ѿ��s��9���Ǿ����P   P   )������.���U������-���I���g��3����������������+���ck���M��m1��9��-��P   P   ٷ���˿�=ҿ��ʿ�&������Ko��^I���&��
��)����辽~澽K꾽�������+���M���s��͘��P   P   ���������������i�������2���̿��f��S	���������Ij���j��҇���������ck��5ѿ�%6��P   P   �i�������4½<O½G3½����e������_%��r�����
����>��(��X@��҇������+����*������P   P   3½d�½�}ý=�ý��ý*{ý��½�.½jP���m�������澽�h��V'��(���j��K꾽���Mr��0U��P   P   �½��ýŪĽH2Ž&`Ž�0ŽǧĽ��ý�½`���_���Ȥ���㾽�h���>��Ij��~澽�������k���P   P   ;=ý
�ĽH�Ž�kƽW�ƽ��ƽ�iƽ��Ž�~Ľ�8ý����X���Ȥ���澽
��������辽���v���Z���P   P   �`ý��Ľ]:ƽ|Rǽ�ȽnGȽBȽ�Oǽ�6ƽY�Ľ�[ý����_������������)�������������P   P   �<ýa�Ľjqƽ��ǽ�Ƚ�TɽATɽ1�Ƚ��ǽ�mƽY�Ľ�8ý`����m��r���S	��
��3���-p�����P   P   [�½,�Ľ�9ƽ��ǽ�ɽ��ɽ�+ʽ{�ɽCɽ��ǽ�6ƽ�~Ľ�½jP��_%���f���&���g��{'��S��P   P   �0½9�ý��ŽJRǽ�Ƚ��ɽzwʽ�vʽ{�ɽ1�Ƚ�Oǽ��Ž��ý�.½�����̿�^I���I���Ϳ�����P   P   Eg����½��Ľxkƽ�Ƚ}UɽI,ʽzwʽ�+ʽATɽBȽ�iƽǧĽ��½�e��2��Ko���-���o���2��P   P   r�������E|ý�1Ž��ƽ>HȽ}Uɽ��ɽ��ɽ�TɽnGȽ��ƽ�0Ž*{ý��������������������P   P   =��������3½��ým`Ž��ƽ�Ƚ�Ƚ�ɽ�Ƚ�ȽW�ƽ&`Ž��ýG3½i���&���U���ľ�k��P   P   ����Cʿ�O����N½��ý�1ŽxkƽJRǽ��ǽ��ǽ|Rǽ�kƽH2Ž=�ý<O½�����ʿ�.���ӈ��ӈ��P   P   +b��^�:ѿ�O����3½E|ý��Ľ��Ž�9ƽkqƽ]:ƽH�ŽŪĽ�}ý�4½����=ҿ�򾽲b��b1��P   P   9���U��^�Cʿ�����������½9�ý,�Ľa�Ľ��Ľ
�Ľ��ýd�½���������˿����V��y��P   P   >���n���S��Q¿��O�����������$½s�½��½�ý��½��½�&½����~���;R��(Ŀ��T��
��P   P   
�����v/���p���˿�;:��ޮ�� ��)���S���9�����������̄��W"��V����<���Ϳ��r���0��P   P   �T��YJ��6T��!q��	����ٿ�G���d��������������	��A�������w���g��c!���ܿ������r��P   P   (Ŀ�پ������¿��˿��ٿ�+뿽~��!���,���<��VE���E��_>���.�������&�ܿ��Ϳ�P   P   ;R���`��|e���_���O���9������ ��翽�ѿ�S���.������p���7ÿ�TԿ�c꿽���c!���<��P   P   ~���� ���:���9��:����������c�����ѿ�����,n���X��&Y���o������TԿ���g��V���P   P   ���������(½<½='½����s����������+��b����m��	9��'���:���o��7ÿ��.��w���W"��P   P   �&½c�½�ý�OýQOý�ý��½(#½���������:�������W���&��'��&Y��p���_>������̄��P   P   ��½�\ý
�ý�XĽ|ĽiWĽ��ý�Yý�½���������B�������W��	9���X������E��A�������P   P   ��½�ý��Ľ�=Ž��Ž��Ž?<ŽͤĽ��ýu�½)���{���B�������m��+n��.���VE���	������P   P   �ýAĽ�Ž��Ž�iƽj�ƽnhƽ��Ž�Ž�Ľ_ý)��������:��b�������S����<������9���P   P   ��½�Ľ�@Ž�>ƽs�ƽ�YǽlYǽ�ƽ�<ƽ�=Ž�Ľu�½��������+��ѿ��ѿ��,������S���P   P   s�½�ýQŽ�>ƽ�)ǽ�ǽ�ǽ=�ǽ(ǽ�<ƽ�Ž��ý�½�����������翽!�����)���P   P   �$½�[ý@�Ľ{�Žx�ƽO�ǽo,Ƚ�+Ƚ=�ǽ�ƽ��ŽͤĽ�Yý(#½����c��� ��~���d�� ��P   P   ����8�½�ýt=Ž�iƽkZǽH�ǽo,Ƚ�ǽlYǽnhƽ?<Ž��ý��½s���������+뿽G��ޮ��P   P   ��������ý�XĽO�Ž�ƽkZǽO�ǽ�ǽ�Yǽj�ƽ��ŽiWĽ�ý���������9���ٿ��ٿ�;:��P   P   �O��z��|'½WOý:|ĽO�Ž�iƽx�ƽ�)ǽs�ƽ�iƽ��Ž|ĽQOý='½:���O���˿�	����˿�P   P   Q¿��_��r9���;½WOý�XĽt=Ž{�Ž�>ƽ�>ƽ��Ž�=Ž�XĽ�Oý<½�9���_���¿�!q���p��P   P   �S�������d��r9��|'½�ý�ý@�ĽQŽ�@Ž�Ž��Ľ
�ý�ý�(½�:��|e�����6T��v/��P   P   n��~I�������_��z�����8�½�[ý�ý�ĽAĽ�ý�\ýc�½����� ���`��پ��YJ�����P   P   쿿�Vҿ����Z������I9������½�u½ȭ½#�½	�½jv½>½s����:��|���s[��W���ҿ�P   P   �ҿ��ҿ��뿽[��Ua���������{]�������������������������/_���
��r����b������쿽P   P   W��< ��������@��7l������������)��2C���K���C���*���������y���tn��B�����P   P   s[��W���V��?Z��a��l���z�����������������	���h�������J���^��������|��tn���b��P   P   |�������1�����������U����������:u��ye���X���Q��>O���R���Z���g���w������y���r���P   P   �:��I]���o��o��&\���8��1�����x���$e��9������
���
�����&;���g��^��������
��P   P   s���o���<½�-½1½�������o\��� ��[���DX�����O�忽�󿽦���Z��J������/_��P   P   >½m�½��½��½��½x�½@�½|½�����'������P���	���俽忽�
���R�������*������P   P   jv½�ýsýܻý��ý��ýpqýj ý�s½�����@��$���PM���	��O򿽥
��>O��h����C������P   P   �½o^ý��ý�cĽ��Ľ �ĽTbĽ`�ý�[ý �½D���LI��$����P���������Q��	����K�����P   P   #�½�ý�HĽ��Ľ�=ŽC^Ž�<Ž�Ľ�FĽs�ý��½D����@�����DX��9���X������2C������P   P   ȭ½��ý�eĽ'ŽG�Ž)�Ž��ŽB�Ž^ŽJcĽs�ý �½�����'��[���$e��ye������)������P   P   �u½�]ý�HĽŽ��Ž�7ƽ{]ƽ�6ƽ��Ž^Ž�FĽ�[ý�s½����� ��x���:u�������������P   P   �½ýM�ýq�Ľ[�Ž�7ƽP�ƽ	�ƽ�6ƽB�Ž�Ľ`�ýj ý|½o\����������������{]��P   P   ���v�½Rrý;cĽ+>Ž��Ž�]ƽP�ƽ{]ƽ��Ž�<ŽTbĽpqý@�½���1������z��������P   P   I9��3���/�½��ýʜĽ�^Ž��Ž�7ƽ�7ƽ)�ŽC^Ž �Ľ��ýx�½�����8��U���l��7l������P   P   ����K\��H½��½��ýʜĽ+>Ž[�Ž��ŽG�Ž�=Ž��Ľ��ý��½1½&\������a��@��Ua��P   P   Z�������n���-½��½��ý;cĽq�ĽŽ'Ž��Ľ�cĽܻý��½�-½o������?Z�����[��P   P   ���)V��r����n��H½/�½RrýM�ý�HĽ�eĽ�HĽ��ýsý��½<½�o��1����V������뿽P   P   Vҿ�~���)V������K\��3���v�½ý�]ý��ý�ýo^ý�ým�½o���I]������W��< ���ҿ�P   P   �W��&e��׋��o���E��o��w���"½�X½`�½��½��½�Y½
½����fp��v��y���z����e��P   P   �e��_e��Ix��<�������M���L��x���3�������n�������0���R���׋��.N���������m���y��P   P   z�������΋������������������"��G���c��"v���|���v���d��rH��v$��������������m���P   P   y���>����������b����������&�����������������������N���!��������������P   P   v��k ��#�������O��������������F���{�������
���Y����������l���!����������P   P   fp������H���Җ��ވ���n���K��I"������ ���������J����������^������N���v$��-N��P   P   ����N����½K$½½������������3F�������������B|��4s���|�����������rH��׋��P   P   
½�d½��½��½[�½z�½�b½�½ǽ��Tb���
�����������r��4s������Y�������d��R���P   P   �Y½��½býUIýZý�Hý'ý��½�W½���yt�������������B|��J���
�������v��0���P   P   ��½&ý�qý2�ý�ý��ý�ý}pý5ý8�½�����z������������������������|������P   P   ��½$'ý¯ý�Ľ�bĽ�{ĽebĽtĽ�ý8%ý��½����yt���
���������{�����"v��n���P   P   `�½�&ý|�ýLĽ��Ľ��Ľ7�ĽҭĽ�JĽ��ý8%ý8�½���Tb����� ���F�������c������P   P   �X½�ý��ý	LĽ\�Ľ�Ž�3Ž;ŽB�Ľ�JĽ�ý5ý�W½ǽ��3F��������������G��3���P   P   "½��½�qý�Ľ��Ľ�ŽWRŽXRŽ;ŽҭĽtĽ}pý��½�½����I"������&����"��x���P   P   w����c½�ý��ýCcĽ��Ľ�4ŽWRŽ�3Ž7�ĽebĽ�ý'ý�b½�����K��������������L��P   P   o��{����½KIýA�ý#|Ľ��Ľ�Ž�Ž��Ľ�{Ľ��ý�Hýz�½�����n��O���������M��P   P   E�����½s�½ZýA�ýCcĽ��Ľ\�Ľ��Ľ�bĽ�ýZý[�½½ވ����b�����������P   P   o����������C$½s�½KIý��ý�Ľ	LĽLĽ�Ľ2�ýUIý��½K$½Җ�������������<���P   P   ׋�������"������½�½�ý�qý��ý|�ý¯ý�qýbý��½�½H���#�����΋��Ix��P   P   &e���������������{����c½��½�ý�&ý$'ý&ý��½�d½N�������k ��>�������_e��P   P   U���G�����������U��/���F����½C½mb½�l½�b½�C½½@���U����V�����#�������P   P   �����������~���9 ��,M��<}����������������������������)���+~���N��{!��Z������P   P   #������������������'��5C���^��_y������������������\z��W`��{D��@(�����Z���P   P   ���u��h�����, ���&��#.��^7��A@���G���M��Q��PQ���N���H���A���8���/��@(��{!��P   P   �V���\��L^��
\���U��PM���B��l7��-��"��B��������-�����#���.���8��{D���N��P   P   U������A�������/��� ����|���^���?��"���
��o���(�������f�������#���A��W`��+~��P   P   @�������}½�½½^�������i����x��!G�����=������5���W���f������H��\z��)���P   P   ½�L½�t½��½%�½�s½dK½v½��� ��� M������������5�������-���N���������P   P   �C½�½z�½t�½ý��½g�½A�½2B½m���r����O������������(������PQ��������P   P   �b½��½�ý�Mý{mýDmý�Lý�ý��½�`½D��������O����=���o������Q��������P   P   �l½��½�?ý�ý�ý�ý��ýюý^>ý^�½Fk½D���r��� M������
��B���M����������P   P   mb½��½vOý�ý��ý� ĽA Ľ:�ýA�ý)Ný^�½�`½m��� ���!G��"��"���G���������P   P   C½��½�?ý%�ýĽ�GĽ�[ĽZGĽĽA�ý^>ý��½2B½����x���?��-��A@��_y������P   P   �½`�½�ýˏý��ý�GĽ�qĽ�qĽZGĽ:�ýюý�ýA�½v½i����^��l7��^7���^������P   P   F����K½$�½eMý%�ý� Ľ�\Ľ�qĽ�[ĽA Ľ��ý�Lýg�½dK½�����|���B��#.��5C��<}��P   P   /�������ft½e�½�mý��ý� Ľ�GĽ�GĽ� Ľ�ýDmý��½�s½^��� ���PM���&��'��,M��P   P   �U��6���½K�½Dý�mý%�ý��ýĽ��ý�ý{mýý%�½½/����U��, �����9 ��P   P   ����[��ҳ���½K�½e�½eMýˏý%�ý�ý�ý�Mýt�½��½�½����
\���������~���P   P   ���� ��/^��ҳ��½gt½$�½�ý�?ývOý�?ý�ýz�½�t½}½A���L^��h����������P   P   G������� ���[��6��������K½`�½��½��½��½��½�½�L½��������\��u���������P   P   ���"���7��Z��������������½@3½�I½�P½�I½�3½½g�������l����Z���8��U"��P   P   U"��N"���+��-@��]\���}�������������-���v ½� ½����]������������~��s]���@��^,��P   P   �8���4��8��)@���N���a��Ov�����D�������ɷ���������Q������1���`w���b���O���@��P   P   �Z���W���W��.Z��s\���a���f��Sm��t��fy��M~��_��������~��Oz��u���n���g���b��s]��P   P   l���2���
������������}��	v��um��]e���^��qY���U���T��V��Z���_��uf���n��`w���~��P   P   ����������������!�������c���ڊ��[s���^��L��P>���8��9��%?���L���_��u��1�������P   P   g�������½�½�½����*���c�������.y���X��8>��L/���)���/��%?��Z��Oz���������P   P   ½:½�W½�h½2h½UW½J9½�½���������}��PU��y8��$)���)��9��V���~��Q���]���P   P   �3½}k½j�½��½Ͼ½K�½i�½$j½[2½C����������S��y8��L/���8���T�������������P   P   �I½�½��½��½;ýý�½N�½Ȏ½sH½>����������PU��8>��P>���U��_�������� ½P   P   �P½r�½��½m'ýQMý�Yý�Lý�&ýe�½e�½�O½>�������}���X��L��qY��M~��ɷ��v ½P   P   �I½��½��½l@ýFvý<�ý�ý�uý�?ý�½e�½sH½C�������.y���^���^��fy������-���P   P   @3½��½Q�½e@ýN�ý��ý��ýB�ý��ý�?ýe�½Ȏ½[2½��������[s��]e��t��D�������P   P   �½�j½��½l'ýuvýv�ý��ý��ýB�ý�uý�&ýN�½$j½�½c���ڊ��um��Sm���������P   P   �����9½)�½��½0Mý[�ý�ý��ý��ý�ý�Lý�½i�½J9½*���c���	v���f��Ov�����P   P   ����9����W½x�½GýZý[�ýv�ý��ý<�ý�YýýK�½UW½���������}���a���a���}��P   P   ���-����½Zh½�½Gý0MýuvýN�ýFvýQMý;ýϾ½2h½�½!�������s\���N��]\��P   P   Z��a���i����½Zh½x�½��½l'ýe@ýl@ým'ý��½��½�h½�½��������.Z��)@��-@��P   P   �7���W�����i����½�W½)�½��½Q�½��½��½��½j�½�W½½����
����W��8���+��P   P   "���4���W��a���-���9����9½�j½��½��½r�½�½}k½:½��������2����W���4��N"��P   P   �W���]���m������B����������½�'½Q8½r>½�8½�'½#½�����������������m���]��P   P   �]���]��;f���t��_�������*���r�������S���|½�½�����������¼���������u���f��P   P   �m���j���m���t��)�����������������$���h���������������!���y���Ҝ��L������u��P   P   ��������v�����������������������������q���n�������ˡ��`�������̖�����L������P   P   ����@���1�������������ۛ������������6����������0���͆��a���܏��̖��Ҝ������P   P   ����A���C���*�������������c���:�������l}���s��?n��Rn��:t��
~��a�������y���¼��P   P   ����� ½�½�½�½8 ½�������;���z��������s���g���b���g��:t��͆��`���!������P   P   #½,½�B½�M½�M½�B½\+½>½]���t���Ҡ�������m��qb���b��Rn��0���ˡ����������P   P   �'½RQ½(r½	�½y�½��½bq½oP½�&½��������Ң������m���g��?n������������������P   P   �8½�l½��½��½Y�½4�½E�½�½�k½�7½�½����Ң�������s���s�����n��������½P   P   r>½�y½ȯ½�½~�½ý%�½��½��½�x½c=½�½����Ҡ������l}��6���q���h���|½P   P   Q8½�y½�½��½TýT(ýB(ý�ý��½j�½�x½�7½����t���z��������������$���S���P   P   �'½<l½ʯ½m�½wýh>ýoIý1>ýý��½��½�k½�&½]���;���:�������������������P   P   �½�P½��½�½_ý�>ýUý�Tý1>ý�ý��½�½oP½>½���c�������������r���P   P   ����+½�q½��½x�½�(ýiIýUýoIýB(ý%�½E�½bq½\+½�������ۛ��������*���P   P   ���x ½�B½׆½r�½+ý�(ý�>ýh>ýT(ýý4�½��½�B½8 ½�������������������P   P   B��������½�M½��½r�½x�½_ýwýTý~�½Y�½y�½�M½�½�����������)��_���P   P   �����������w½�M½׆½��½�½m�½��½�½��½
�½�M½�½*�����������t���t��P   P   �m��@���"�������½�B½�q½��½ʯ½�½ȯ½��½(r½�B½�½C���1���v����m��;f��P   P   �]���j��@�����������x ½�+½�P½<l½�y½�y½�l½RQ½,½� ½A���@��������j���]��P   P   ����������0���d���k���n����½�½�*½b/½�*½�½�½���������������r���	���P   P   	����������̚��R���&�������/�������x����½ ½������������R������������������P   P   r�������I�������k�����������$�������X����������,�������C����������D���0������P   P   ����=������4���i�������,��������������p���_�����������|�������1������D�������P   P   ���@���J������j����������x���1����������V���������������A���	���1����������P   P   ���� ���E��� �������?�������������������������ߕ��ܕ��O���$���A�����������R���P   P   ����5½�½�½c½�½�������]�������ȧ������e���5������O�������|���C�������P   P   �½�"½_2½�:½�:½2½"½�½>�����������������@���5���ܕ������������������P   P   �½F=½xU½�e½�k½:e½U½�<½½����V�������������e���ߕ����������,�������P   P   �*½�P½]q½��½!�½�½=�½�p½P½M*½V½R����������������V���_������ ½P   P   b/½C[½ك½O�½b�½Y�½/�½��½U�½�Z½q.½V½V������ȧ���������p��������½P   P   �*½[½O�½�½]�½��½��½��½V�½ƈ½�Z½M*½�����������������������X���x���P   P   �½�P½��½԰½a�½q�½��½Y�½8�½V�½U�½P½½>���]������1���������������P   P   �½4=½#q½E�½B�½��½0�½ �½Y�½��½��½�p½�<½�½��������x�������$���/���P   P   n���|"½QU½��½��½�½y�½0�½��½��½/�½=�½U½"½�����������,�����������P   P   k����½<2½|e½H�½E�½�½��½q�½��½Y�½�½:e½2½�½?��������������&���P   P   d��������½�:½�k½H�½��½B�½a�½]�½b�½!�½�k½�:½c½����j���i���k���R���P   P   0����������½�:½|e½��½E�½԰½�½O�½��½�e½�:½�½ ������4�������̚��P   P   ��� ����������½<2½QU½#q½��½O�½ك½]q½xU½_2½�½E���J������I�������P   P   ������� �����������½|"½4=½�P½[½C[½�P½F=½�"½5½ ���@���=����������P   P   ��������������k������������	½�½�!½�$½�!½)½q
½������������q���S���ڪ��P   P   ڪ���������c���A���w�����������m�������½1½
 ½d�����������������������)���P   P   S������F���C���b�����������p�������9�������-������������������8���	����������P   P   q���ɿ���������@����������� ��������������������������l������v���f���	�������P   P   ��������\�����������%���������������������U�����������������������v���8�������P   P   ��������������������C��������������A�������b���U���Y���k���@������������������P   P   �����½p
½7½H
½�½����<�����������$���(���(�����������k�������l�����������P   P   q
½l½f&½�-½s-½&½�½�	½������P������
���ۭ������Y���������������d���P   P   )½/½HA½HL½P½�K½A½�.½`½H���a���Y���|���
���(���U��������������
 ½P   P   �!½W=½�U½g½zo½wo½�f½�T½�<½-!½�½����Y������(���b���U�������-���1½P   P   �$½�E½�b½�y½ǈ½��½��½by½-b½)E½8$½�½a���P���$������������������½P   P   �!½�E½#g½s�½W�½��½��½ �½�½�f½)E½-!½H����������A����������9�������P   P   �½M=½�b½��½˞½��½��½�½��½�½-b½�<½`½����������������������m���P   P   �	½)/½sU½�y½-�½��½q�½@�½�½ �½by½�T½�.½�	½<���������� ���p�������P   P   ����5½A½
g½ֈ½�½�½q�½��½��½��½�f½A½�½������������������������P   P   �����½I&½AL½�o½�½�½��½��½��½��½wo½�K½&½�½C���%�����������w���P   P   k�������e
½�-½�O½�o½ֈ½-�½˞½W�½ǈ½zo½P½s-½H
½��������@���b���A���P   P   �����������½�-½AL½
g½�y½��½s�½�y½g½HL½�-½7½�����������C���c���P   P   ���������������e
½I&½A½sU½�b½#g½�b½�U½HA½f&½p
½����\�������F������P   P   ����	����������������½5½)/½M=½�E½�E½W=½/½l½�½��������ɿ���������P   P   ���������������������������	½�½i½�½}½L½�	½���/������^����������P   P   ����x�������A���4���]���O������������½ ½1½�½���������������}�����������P   P   ����������C�������������������&�������.���(���K���
����������a���;���$�������P   P   ^��������������#�����������!�������W������� ���'�����������c���}�������;���}���P   P   ����������������������������������������������>���D����������}���a�������P   P   /���������������(�������x���}���<�������a������������������������c����������P   P   ���d½S	½�
½O	½)½���������������������������O����������D��������������P   P   �	½�½V½Y#½)#½½s½g	½9�������r�������x���r���O�������>�������
�������P   P   L½q$½u1½:½<½�9½,1½8$½�½½������������x���������������'���K����½P   P   }½</½�@½FM½�T½|T½M½;@½�.½½�½���������������������� ���(���1½P   P   �½Z4½UJ½B[½�f½#k½�f½#[½J½�3½L½�½����r������a�����������.��� ½P   P   i½Z4½�M½�c½�r½Qz½bz½Kr½Cc½RM½�3½½½����������������W��������½P   P   �½G/½*J½�c½�v½��½��½~�½�v½Cc½J½�.½�½9�������<����������&�������P   P   �	½y$½�@½q[½mr½��½��½b�½~�½Kr½#[½;@½8$½g	½����}�������!�����������P   P   �����½D1½[M½�f½�z½��½��½��½bz½�f½M½,1½s½����x���������������O���P   P   ���½5½:½�T½Ok½�z½��½��½Qz½#k½|T½�9½½)½���������������]���P   P   ����&���i	½@#½<½�T½�f½mr½�v½�r½�f½�T½<½)#½O	½(������#�������4���P   P   ������������
½@#½:½[M½q[½�c½�c½B[½FM½:½Y#½�
½�����������C���A���P   P   ����������������i	½5½D1½�@½*J½�M½UJ½�@½u1½V½S	½������������������P   P   ����������������&���½�½y$½G/½Z4½Z4½</½q$½�½d½����������������x���P   P   ~�����������7����������������	½=½w½B½�½G½�	½�����������a����������P   P   ����������������Z���H�������f���(���X½�½�½i½t�����������h�������?�������P   P   �����������	���%�������}����������������������������������� �������P���!���?���P   P   a�����������<���K�������5�����������@���������������1���x���F�������J���P�������P   P   ����
��������������"�������l���������������{���9���u�����������-�����������h���P   P   ���������������h�������������������p������>���O�������l���d�������F��� �������P   P   �����½d	½�	½N	½�½d���=�������	�������;�������U�������l�������x�����������P   P   �	½�½�½7½	½~½l½�	½���r����������6���G���U�������u���1�������t���P   P   G½�½c&½�,½c/½�,½
&½�½�½½����v���T���6�������O���9�����������i½P   P   �½�$½�1½�:½�?½�?½�:½�1½�$½c½�½����v������;���>���{������������½P   P   B½1)½�8½�E½8M½qO½%M½�E½�8½�(½�½�½����������������������������½P   P   w½K)½B;½�J½1V½X\½e\½�U½GJ½;½�(½c½½r���	���p�������@�������X½P   P   =½�$½�8½{J½�X½�b½1f½�b½�X½GJ½�8½�$½�½�����������������������(���P   P   �	½�½�1½�E½2V½�b½�g½�g½�b½�U½�E½�1½�½�	½=�������l�����������f���P   P   �����½V&½�:½M½o\½f½�g½1f½e\½%M½�:½
&½l½d�����������5���}�������P   P   �����½�½�,½�?½�O½o\½�b½�b½X\½qO½�?½�,½~½�½����"�����������H���P   P   ����j���b	½(½�/½�?½M½2V½�X½1V½8M½�?½c/½	½N	½h�������K���%���Z���P   P   7������������	½(½�,½�:½�E½{J½�J½�E½�:½�,½7½�	½��������<���	�������P   P   ����������������b	½�½V&½�1½�8½B;½�8½�1½c&½�½d	½�������������������P   P   ����s�����������j����½�½�½�$½K)½1)½�$½�½�½�½����
���������������P   P   L���.�������1���(��������½�½g½�½�½½I½o½�½���.���F�������:���P   P   :���3������x�����������Z���3���½�½!½�½�½�½g���u���%����������+���P   P   ������������~���o���Q���g���r�����������j�������������������������������y�������P   P   F������o���<�������K���
���@���"���~�������|���������������s�������/����������P   P   .������>��������������X���E����������������� �����������-���(�����������%���P   P   ���P���k�������$�������I���_��������������������O���P��� ���-���s�������u���P   P   �½�½�½
½�½�½�½�������q���z������������������P���������������g���P   P   o½�½½#½
½�½�½L½½~����������� �����������O����������������½P   P   I½b½�½j"½�$½�"½�½½½]½L���/���6��� ����������� ������������½P   P   ½�½Q&½�-½e1½1½{-½H&½�½�½�½s���/����������������|��������½P   P   �½' ½2+½65½o;½h=½�;½5½�*½�½H½�½L�������z��������������j���!½P   P   �½6 ½�-½t9½�A½�E½�E½KA½.9½�-½�½�½]½~���q�����������~��������½P   P   g½�½8+½P9½�C½�J½8L½�J½D½.9½�*½�½½½����������"�������½P   P   �½½3&½<5½�A½�J½�O½�O½�J½KA½5½H&½½L½���_���E���@���r���3���P   P   �½�½½�-½t;½�E½OL½�O½8L½�E½�;½{-½�½�½�½I���X���
���g���Z���P   P   �����½�½R"½?1½�=½�E½�J½�J½�E½h=½1½�"½�½�½��������K���Q�������P   P   (���0����½(½�$½?1½t;½�A½�C½�A½o;½e1½�$½
½�½$����������o�������P   P   1�������u���
½(½R"½�-½<5½P9½t9½65½�-½j"½#½
½��������<���~���x���P   P   ����i���F���u����½�½½3&½8+½�-½2+½Q&½�½½�½k���>���o����������P   P   .�������i�������0����½�½½�½6 ½' ½�½b½�½�½P�������������3���P   P   ����������������������[½D½%½G½�½j½½%½s½!�����������C�������P   P   ����������������f������x���)���½�½�½�½ ½S½Q�������E���������������P   P   C���F���1������������������L���$����������c���:�������5���������������������P   P   ����s���l�������s�����������X������O�����������������������*������������������P   P   ��������������������"�������i������������������������&���K��������������E���P   P   !���0������������������T���i����������a���2���.���e�������Z���K���*�����������P   P   s½½W½]	½J½
½L½�������]�������K���Q���,����������&�������5���Q���P   P   %½�½1½7½ ½�½A½½½������������7�������,���e���������������S½P   P   ½'½4½�½d½½0½�½�½�½����W�������7���Q���.�����������:��� ½P   P   j½½�½�#½)&½�%½Z#½y½�½F½{½P���W�������K���2����������c����½P   P   �½�½�"½)½9-½P/½s-½�(½�"½}½x½{½������������a��������������½P   P   G½�½�#½�,½2½"6½�5½�1½d,½�#½}½F½�½����]���������O��������½P   P   %½½�"½�,½�3½�8½O:½�8½�3½d,½�"½�½�½½���������������$���½P   P   D½�½½)½$2½�8½�<½=½�8½�1½�(½y½�½½���i���i���X���L���)���P   P   [½8½v½�#½l-½�5½�:½�<½O:½�5½s-½Z#½0½A½L½T��������������x���P   P   ����(½½�½&½m/½�5½�8½�8½"6½P/½�%½½�½
½����"��������������P   P   ������1½/½�½&½l-½$2½�3½2½9-½)&½d½ ½J½�������s�������f���P   P   ������������e	½/½�½�#½)½�,½�,½)½�#½�½7½]	½��������������������P   P   ���f�����������1½½v½½�"½�#½�"½�½4½1½W½��������l���1�������P   P   ����K���f����������(½8½�½½�½�½½'½�½½0�������s���F�������P   P   1���y�����������B���$ ½t½<	½d½'½�½½}½?	½�½U ½3������ ���~���P   P   ~���u���U�����������������D½½½]½s½F½
½[½���!�����������b���P   P    ���Q���������������w������9���y�������� ½T ½� ½��������x���=��������������P   P   �������������������y���p���m�������K����������������������������������������P   P   3���������������:���������l�������1����������������������k�����������=���!���P   P   U ½�½�½�½�½/ ½����\�������b�����������#���&���$�������k�������x������P   P   �½�½s½�½�½�½s½1½U���V���V�������&����������$��������������[½P   P   ?	½�½�½�½�½z½�½	½�½������������#�����������&��������������
½P   P   }½�½½�½½�½½�½?½½� ½��������#���&���#����������� ½F½P   P   ½1½�½�½�½�½�½�½½�½J½, ½�����������������������T ½s½P   P   �½½�½� ½�#½>$½�#½� ½�½�½h½J½� ½����V���������������� ½]½P   P   '½�½1½8"½�'½�)½�)½�'½/"½½�½�½½����V���b���1���K�������½P   P   d½/½�½U"½�(½�,½v-½�,½n(½/"½�½½?½�½U���������������y���½P   P   <	½�½�½� ½�'½�,½.½.½�,½�'½� ½�½�½	½1½\���l���m���9���D½P   P   t½�½½�½�#½�)½�-½.½v-½�)½�#½�½½�½s½�������p���������P   P   $ ½�½�½�½�½,$½�)½�,½�,½�)½>$½�½�½z½�½/ ½���y���w������P   P   B����½n½�½;½�½�#½�'½�(½�'½�#½�½½�½�½�½:���������������P   P   ���������½	½�½�½�½� ½U"½8"½� ½�½�½�½�½�½����������������P   P   �������������½n½�½½�½�½1½�½�½½�½s½�½������������U���P   P   y���Y������������½�½�½�½/½�½½1½�½�½�½�½��������Q���u���P   P   h�����������m���H����½�½L½�
½�½½i½�
½s½�½�½e���������������P   P   ��������(����������4���+½W½½f½ ½c½�½�½[½!½F����������N���P   P   ���������������?���t���}�������J½X½�½�½�½d½�½ ½��������W������P   P   ����;��� ���j�������l�������F���z���M�������������������g���f���M���������������P   P   e���s��� ½����S���2�������5����������������������������������B���M�������F���P   P   �½�½�½�½�½�½
½����a�������*���q���}���Q���o���d�������f��� ½!½P   P   �½�½�½�½�½�½�½M½B½<�������^����������K���o�������g����½[½P   P   s½c½e½U½\½c½]½F½�½`½b�������k�����������Q����������d½�½P   P   �
½w½u½�½T½�½S½j½�
½U½�½����@���k������}������������½�½P   P   i½�½'½�½½.½�½�½�½`½6½m½��������^���q������������½c½P   P   ½m½q½½½�½�½½c½1½�½6½�½b�������*������������½ ½P   P   �½8½�½&½F½Z ½o ½a½½�½1½`½U½`½<�����������M���X½f½P   P   �
½q½�½B½% ½x"½
$½w"½�½½c½�½�
½�½B½a�������z���J½½P   P   L½�½?½�½3½�"½f%½B%½w"½a½½�½j½F½M½����5���F�������W½P   P   �½~½3½�½½� ½�#½f%½
$½o ½�½�½S½]½�½
½��������}���+½P   P   �½�½f½�½½�½� ½�"½x"½Z ½�½.½�½c½�½�½2���l���t���4���P   P   H����½�½E½F½½½3½% ½F½½½T½\½�½�½S�������?�������P   P   m��������½�½E½�½�½�½B½&½½�½�½U½�½�½����j���������P   P   ������� ½�½�½f½3½?½�½�½q½'½u½e½�½�½ ½ �������(���P   P   ����������������½�½~½�½q½8½m½�½w½c½�½�½s���;�����������P   P   ��������6�������v½P½�½b½?
½�½�½�½c
½�½�½H½�½ ½�������P   P   ������������h���� ½�½{½d½�½�½i½�½�½�½f½�½�½} ½��������P   P   �������������� ½ ½x½>½-½�½B½�½+½�½N½M½�½) ½Y ½����P   P    ½�������� ½� ½ ½� ½3½½�½!½�½�½&½½*½D½� ½) ½} ½P   P   �½-½½>½m½�½�½)½½� ½���� ½����F ½����� ½)½D½�½�½P   P   H½�½}½l½�½M½_½3½½� ½R�����������l������������ ½*½M½�½P   P   �½�½u½�½>½�½�½e½5½[½�������� �������[�����������½N½f½P   P   �½'
½�½�½½�½)
½s½�½�½�½ ½�����������l���F ½&½�½�½P   P   c
½�½[½t½e½2½7½�½[
½�½#½�½�������� ������������½+½�½P   P   �½�½½[½�½�½�½�½�½�½�½e½�½ ½�������� ½�½�½�½P   P   �½d½�½�½�½"½b½�½�½<½�½�½#½�½����R�������!½B½i½P   P   �½A½�½�½C½�½�½I½�½�½<½�½�½�½[½� ½� ½�½�½�½P   P   ?
½�½�½�½�½½½½�½�½�½�½[
½�½5½½½½-½�½P   P   b½�½5½�½;½½�½�½½I½�½�½�½s½e½3½)½3½>½d½P   P   �½O
½½Y½�½½�½�½½�½b½�½7½)
½�½_½�½� ½x½{½P   P   P½�½�½�½	½�½½½½�½"½�½2½�½�½M½�½ ½ ½�½P   P   v½�½M½�½½	½�½;½�½C½�½�½e½½>½�½m½� ½ ½� ½P   P   ����@½X½�½�½�½Y½�½�½�½�½[½t½�½�½l½>½ ½����h���P   P   6�������-½X½M½�½½5½�½�½�½½[½�½u½}½½�����������P   P   ����e�������@½�½�½O
½�½�½A½d½�½�½'
½�½�½-½������������P   P   ���^ ½^½�½�½2½;½�½�	½�
½�½�
½�	½�½=½+½�½�½J½] ½P   P   ] ½| ½� ½�½(½�½½�½d½�½½�½�½b½�½½�½�½�½½P   P   J½E½/½�½�½�½�½I½�½Z½�½*½�½�½�½G½�½�½�½�½P   P   �½½½�½	½�½�½�½�½M½2½�½�½&½C½�½�½½�½�½P   P   �½"½�½%½�½�½�½�½�½=½�½�½{½�½�½I½p½�½�½�½P   P   +½�½�½�½½2½�½D½�½*½�½�½�½�½�½�½I½�½G½½P   P   =½�½h	½�½9	½�½3½�½�½4½�½�½� ½{ ½� ½�½�½C½�½�½P   P   �½�
½i½½S½l½�
½�½"½�½½�½�½� ½{ ½�½�½&½�½b½P   P   �	½½^½�½�½�½b½�½
½�½�½�½i½�½� ½�½{½�½�½�½P   P   �
½�½�½�½�½�½ ½�½�½m
½�½½�½�½�½�½�½�½*½�½P   P   �½�½�½b½�½�½�½9½�½�½�½�½�½½�½�½�½2½�½½P   P   �
½�½S½-½�½�½�½�½.½-½�½m
½�½�½4½*½=½M½Z½�½P   P   �	½�½�½+½�½p½i½f½�½.½�½�½
½"½�½�½�½�½�½d½P   P   �½½½N½�½V½-½8½f½�½9½�½�½�½�½D½�½�½I½�½P   P   ;½�
½2½�½�½�½�½-½i½�½�½ ½b½�
½3½�½�½�½�½½P   P   2½�½g½�½�½�½�½V½p½�½�½�½�½l½�½2½�½�½�½�½P   P   �½½B	½@½�½�½�½�½�½�½�½�½�½S½9	½½�½	½�½(½P   P   �½!½�½�½@½�½�½N½+½-½b½�½�½½�½�½%½�½�½�½P   P   ^½½�½�½B	½g½2½½�½S½�½�½^½i½h	½�½�½½/½� ½P   P   ^ ½5½½!½½�½�
½½�½�½�½�½½�
½�½�½"½½E½| ½P   P   �½�½*½ ½�½½�½�½�	½-
½�	½e
½�	½�½�½½�½)½F½�½P   P   �½�½�½�½D½�½'½�½u½�½�½�½�½�½½.½�½E½�½�½P   P   F½½½�½-½�½�½p½&½½�½[½�½M½�½p½�½�½C½�½P   P   )½s½�½+½4½�½�½�½�½|½1½t½½#½{½�½½�½�½E½P   P   �½v½�½h½p½�½y½�½�½3½�½�½�½�½�½L½�½½�½�½P   P   ½�½�½e½�½½	½|½�½7½½½�½�½�½½L½�½p½.½P   P   �½e½�½	½	½D½�½�½	½�½�½�½�½�½�½�½�½{½�½½P   P   �½�	½�
½�½�½�
½�	½�½T½+½½�½�½�½�½�½�½#½M½�½P   P   �	½�½6½)½,½½R½�½�	½�½�½n½�½�½�½�½�½½�½�½P   P   e
½�½]½�½O½\½�½f½�½
½�½f½n½�½�½½�½t½[½�½P   P   �	½�½�½$½½�½½�½�½�½�	½�½�½½�½½�½1½�½�½P   P   -
½ ½�½�½½�½�½8½�½�½�½
½�½+½�½7½3½|½½�½P   P   �	½�½�½�½�½½�½½G½�½�½�½�	½T½	½�½�½�½&½u½P   P   �½�½z½(½B½�½�½�½½8½�½f½�½�½�½|½�½�½p½�½P   P   �½�	½?½�½�½�½�½�½�½�½½�½R½�	½�½	½y½�½�½'½P   P   ½L½�
½)½R½�½�½�½½�½�½\½½�
½D½½�½�½�½�½P   P   �½�½ 	½�½/½R½�½B½�½½½O½,½�½	½�½p½4½-½D½P   P    ½i½z½	½�½)½�½(½�½�½$½�½)½�½	½e½h½+½�½�½P   P   *½�½�½z½ 	½�
½?½z½�½�½�½]½6½�
½�½�½�½�½½�½P   P   �½½�½i½�½L½�	½�½�½ ½�½�½�½�	½e½�½v½s½½�½P   P   �½l½[½�½�½'½�½4	½�	½+
½�
½�
½j	½	½�½;½`½�½z½p½P   P   p½l½�½'½�½½ ½r½�½y½�½�½Z½�½�½½½½(½�½P   P   z½½d½&½L½�½½�½½8½{½½�½T½�½�½!½y½6½'½P   P   �½K½k½�½�½q½�½Z½\½�½½1½M½�½�½�½b½�½y½½P   P   `½�½�½z½�½½½e½�½�½<½½�½�½T½�½�½b½!½½P   P   ;½½E½:½½$½	½�½7½�½�½�½½½�½�½�½�½�½½P   P   �½�½�½e	½	½�½�½�½�½½½�½8½�½½�½T½�½�½�½P   P   	½�	½^
½ ½�
½R
½ 
½	½�½½½½½�½�½½�½�½T½�½P   P   j	½�
½½S½9½V½½�
½�	½�½v½.½v½½8½½�½M½�½Z½P   P   �
½n½�½�½�½�½�½�½i½)
½�½!½.½½�½�½½1½½�½P   P   �
½�½�½�½�½F½w½�½�½½�
½�½v½½½�½<½½{½�½P   P   +
½7½�½�½�½�½�½�½�½�½½)
½�½½½�½�½�½8½y½P   P   �	½�½�½�½R½%½[½½	½�½�½i½�	½�½�½7½�½\½½�½P   P   4	½�
½�½�½�½�½½/½½�½�½�½�
½	½�½�½e½Z½�½r½P   P   �½�	½)½�½l½�½�½½[½�½w½�½½ 
½�½	½½�½½ ½P   P   '½�½_
½2½�½}½�½�½%½�½F½�½V½R
½�½$½½q½�½½P   P   �½�½	½�
½½�½l½�½R½�½�½�½9½�
½	½½�½�½L½�½P   P   �½}½D½\	½�
½2½�½�½�½�½�½�½S½ ½e	½:½z½�½&½'½P   P   [½Y½�½D½	½_
½)½�½�½�½�½�½½^
½�½E½�½k½d½�½P   P   l½½Y½}½�½�½�	½�
½�½7½�½n½�
½�	½�½½�½K½½l½P   P   �½½d½�½^½�½�½U	½X
½F
½�
½�
½>
½F	½�½�½@½�½h½"½P   P   "½½I½6½½n½�½\½b½�½�½�½�½�½^½�½~½7½7½L½P   P   h½F½v½'½�½)½�½�½�½�½R½ ½s½�½�½�½�½½�½7½P   P   �½�½�½�½)½½�½�½k½N½E½#½8½/½K½u½�½�½½7½P   P   @½`½½K½W½j½½�½½A½c½�½s½�½�½Y½½�½�½~½P   P   �½O½>½Y½B½�½�½�½F½[½�½�½o½�½�½l½Y½u½�½�½P   P   �½�	½6	½	½0	½u	½�½H½�½a½F½�½"½�½
½�½�½K½�½^½P   P   F	½,
½�
½t
½U
½�
½/
½<	½y½v½G½�½w½�½�½�½�½/½�½�½P   P   >
½�
½�
½g½�½l½�
½{
½E
½�½h½½b½w½"½o½s½8½s½�½P   P   �
½½�½U½3½B½K½�½½[
½�½½½�½�½�½�½#½ ½�½P   P   �
½½�½#½�½½�½"½Y½(½�
½�½h½G½F½�½c½E½R½�½P   P   F
½,½�½�½�½L½L½½�½�½(½[
½�½v½a½[½A½N½�½�½P   P   X
½%½|½�½�½D½�½@½�½�½Y½½E
½y½�½F½½k½�½b½P   P   U	½k
½�½.½½7½�½�½@½½"½�½{
½<	½H½�½�½�½�½\½P   P   �½
½�
½f½�½K½�½�½�½L½�½K½�
½/
½�½�½½�½�½�½P   P   �½�	½�
½?½0½2½K½7½D½L½½B½l½�
½u	½�½j½½)½n½P   P   ^½?½:	½_
½�½0½�½½�½�½�½3½�½U
½0	½B½W½)½�½½P   P   �½D½E½	½_
½?½f½.½�½�½#½U½g½t
½	½Y½K½�½'½6½P   P   d½�½3½E½:	½�
½�
½�½|½�½�½�½�
½�
½6	½>½½�½v½I½P   P   ½S½�½D½?½�	½
½k
½%½,½½½�
½,
½�	½O½`½�½F½½P   P   }½½�½�½B½	½`	½�	½ 
½
½:
½
½
½

½^	½		½D½�½�½	½P   P   	½½7½�½Q½�½�½	½�½	½�	½�	½)	½�½�½�½�½U½�½;½P   P   �½�½�½t½�½�½�½½e½(½�½S½�½½�½%½d½�½�½�½P   P   �½ ½½�½p½�½�½�½V½�½½i½h½½�½<½�½�½�½U½P   P   D½\½F½Q½,½�½{½�½�½,½f½�½�½�½�½+½�½�½d½�½P   P   		½�½�½�½�½	½�½½K½ ½½~½
½½u½�½+½<½%½�½P   P   ^	½�½�	½
½e	½�½U	½�½�½�½y½r½�½�½�½u½�½�½�½�½P   P   

½�	½9
½�
½�
½]
½	½�	½�½
½½½
½�½�½½�½½½�½P   P   
½e
½½\½T½]½�
½�
½�	½
	½�½_½�½
½�½
½�½h½�½)	½P   P   
½�
½�½�½�½�½�½�½�
½/
½�	½:½_½½r½~½�½i½S½�	½P   P   :
½�
½�½
½9½�½>½*½�½|
½
½�	½�½½y½½f½½�½�	½P   P   
½q
½�½;½�½�½�½�½,½½|
½/
½
	½
½�½ ½,½�½(½	½P   P    
½�
½�½<½n½�½�½�½�½,½�½�
½�	½�½�½K½�½V½e½�½P   P   �	½
½�½½�½�½.½½�½�½*½�½�
½�	½�½½�½�½½	½P   P   `	½	½½�½;½�½�½.½�½�½>½�½�
½	½U	½�½{½�½�½�½P   P   	½�½C
½I½�½�½�½�½�½�½�½�½]½]
½�½	½�½�½�½�½P   P   B½�½t	½�
½L½�½;½�½n½�½9½�½T½�
½e	½�½,½p½�½Q½P   P   �½B½�½
½�
½I½�½½<½;½
½�½\½�
½
½�½Q½�½t½�½P   P   �½½d½�½t	½C
½½�½�½�½�½�½½9
½�	½�½F½½�½7½P   P   ½�½½B½�½�½	½
½�
½q
½�
½�
½e
½�	½�½�½\½ ½�½½P   P   ½�½'½Y½�½�½	½q	½_	½
½+
½�	½�	½�	½ 	½�½�½V½O½�½P   P   �½�½:½q½e½�½�½~	½�	½
½�	½�	½$
½}	½_	½�½�½]½_½#½P   P   O½�½>½J½�½�½�½�½�½�½�½�½�½�½�½�½v½�½½_½P   P   V½�½�½c½x½�½7	½�½6½�½�½x½j½�½�½½�½S	½�½]½P   P   �½½O½z½�½�½�½�½�½�½�½½E½½�½i½�½�½v½�½P   P   �½7	½C	½G	½8	½�½�½�½R½\½½½l½k½�½R½i½½�½�½P   P    	½�	½�	½�	½�	½�	½�½j	½�½�½�½�½½�½.½�½�½�½�½_	½P   P   �	½>
½W
½�	½�	½X
½.
½�	½�	½�½�½�½a½�½�½k½½�½�½}	½P   P   �	½�	½�
½�
½>½�
½�
½$
½C	½�	½�½o½^½a½½l½E½i½�½$
½P   P   �	½�
½+½X½�½�½[½�
½�
½5
½�	½�½o½�½�½½½x½�½�	½P   P   +
½�½�½`½�½�½�½�½�½}½�	½�	½�½�½�½½�½�½�½�	½P   P   
½y½1½/½?½A½^½�½½X½}½5
½�	½�½�½\½�½�½�½
½P   P   _	½�
½�½:½�½*½�½C½½½�½�
½C	½�	½�½R½�½6½�½�	½P   P   q	½/
½ ½z½½l½�½�½C½�½�½�
½$
½�	½j	½�½�½�½�½~	½P   P   	½@
½�
½b½�½j½[½�½�½^½�½[½�
½.
½�½�½�½7	½�½�½P   P   �½�	½Z
½�
½�½�½j½l½*½A½�½�½�
½X
½�	½�½�½�½�½�½P   P   �½5	½�	½�	½½�½�½½�½?½�½�½>½�	½�	½8	½�½x½�½e½P   P   Y½½U	½o	½�	½�
½b½z½:½/½`½X½�
½�	½�	½G	½z½c½J½q½P   P   '½�½4½U	½�	½Z
½�
½ ½�½1½�½+½�
½W
½�	½C	½O½�½>½:½P   P   �½�½�½½5	½�	½@
½/
½�
½y½�½�
½�	½>
½�	½7	½½�½�½�½P   P   �½�½v½	½�½Y	½�	½�	½o
½'
½�	½�	½�
½�	½	½E	½�½	½�½�½P   P   �½�½"½�½$	½r	½J	½	½�	½�	½w	½�	½�	½V	½	½o	½Q	½*	½x½�½P   P   �½�½�½g½}½�½�½�	½I	½b	½M	½�	½.	½O	½r	½�	½	½�½|½x½P   P   	½�½�½�½$	½�½ ½�½�½	½�½F	½<	½	½2	½�½�½�½�½*	½P   P   �½o	½�	½k	½�½?	½�½�½�½B	½�½�½�½�½u½	½6	½�½	½Q	½P   P   E	½d	½I	½<	½K	½=	½z	½�	½�½	½½�½�½�½�½b½	½�½�	½o	½P   P   	½%
½�	½	
½�	½2
½u	½	½0	½	½�½�½	½½	½�½u½2	½r	½	½P   P   �	½r
½
½�
½�
½�	½m
½�	½�	½~	½�½�½�½3½½�½�½	½O	½V	½P   P   �
½�
½\
½�
½½�
½d
½�
½e
½�	½<	½A	½�½�½	½�½�½<	½.	½�	½P   P   �	½�
½�
½
½4½&½½�
½�
½(
½�	½�	½A	½�½�½�½�½F	½�	½�	½P   P   �	½�
½�
½�½�½(½�½½½~
½�	½�	½<	½�½�½½�½�½M	½w	½P   P   '
½�
½O
½�½�½�½½o½�½`
½~
½(
½�	½~	½	½	½B	½	½b	½�	½P   P   o
½�
½½�½�½m½�½½½�½½�
½e
½�	½0	½�½�½�½I	½�	½P   P   �	½�
½�
½�½l½�½½�½½o½½�
½�
½�	½	½�	½�½�½�	½	½P   P   �	½�
½A
½½�½½|½½�½½�½½d
½m
½u	½z	½�½ ½�½J	½P   P   Y	½
½
½�
½3½½½�½m½�½(½&½�
½�	½2
½=	½?	½�½�½r	½P   P   �½F	½�	½�
½�
½3½�½l½�½�½�½4½½�
½�	½K	½�½$	½}½$	½P   P   	½�	½^	½�	½�
½�
½½�½�½�½�½
½�
½�
½	
½<	½k	½�½g½�½P   P   v½�½�	½^	½�	½
½A
½�
½½O
½�
½�
½\
½
½�	½I	½�	½�½�½"½P   P   �½�½�½�	½F	½
½�
½�
½�
½�
½�
½�
½�
½r
½%
½d	½o	½�½�½�½P   P   y	½�½Z	½	½G	½�	½X
½'
½'
½j
½�
½[
½
½0
½\
½�	½Y	½	½_	½�½P   P   �½�½�	½~	½(	½B	½O	½�	½�	½�	½T
½[
½�	½�	½�	½^	½	½6	½�	½~	½P   P   _	½�½v	½�	½�	½p	½O	½�	½�	½�	½�	½	½�	½�	½�	½�	½x	½�	½�	½�	½P   P   	½*	½-	½�½	½�	½
½�	½?	½7	½t	½S	½S	½�	½;	½V	½�	½�	½�	½6	½P   P   Y	½�	½j	½�	½�	½	½i	½�	½4	½R	½3	½�	½P	½�	½/	½7	½E	½�	½x	½	½P   P   �	½�	½�	½�	½�	½�	½o	½�	½r	½5	½�	½q	½�½�½g	½�	½7	½V	½�	½^	½P   P   \
½�	½�	½U
½�	½�	½c
½�	½�	½	½F	½r	½�½�	½�½g	½/	½;	½�	½�	½P   P   0
½�	½7
½h
½O
½
½�	½
½�	½�	½�	½�	½�½�	½�	½�½�	½�	½�	½�	½P   P   
½)
½�
½0½V
½V½�
½:
½)
½�	½�	½K	½c	½�½�½�½P	½S	½�	½�	½P   P   [
½a
½�
½#½�
½�
½½�
½M
½d
½P
½�	½K	½�	½r	½q	½�	½S	½	½[
½P   P   �
½�
½�
½½+½U½;½½½�
½	½P
½�	½�	½F	½�	½3	½t	½�	½T
½P   P   j
½�
½½G½�½w½�½g½*½�½�
½d
½�	½�	½	½5	½R	½7	½�	½�	½P   P   '
½W
½�
½=½�
½½�
½½(½*½½M
½)
½�	½�	½r	½4	½?	½�	½�	½P   P   '
½+
½�
½½t½+½�½�½½g½½�
½:
½
½�	½�	½�	½�	½�	½�	½P   P   X
½�	½�
½(½+½{½�
½�½�
½�½;½½�
½�	½c
½o	½i	½
½O	½O	½P   P   �	½�	½ 
½;½�
½d½{½+½½w½U½�
½V½
½�	½�	½	½�	½p	½B	½P   P   G	½�	½�	½b
½_
½�
½+½t½�
½�½+½�
½V
½O
½�	½�	½�	½	½�	½(	½P   P   	½�	½�	½9
½b
½;½(½½=½G½½#½0½h
½U
½�	½�	½�½�	½~	½P   P   Z	½:	½,	½�	½�	½ 
½�
½�
½�
½½�
½�
½�
½7
½�	½�	½j	½-	½v	½�	½P   P   �½�½:	½�	½�	½�	½�	½+
½W
½�
½�
½a
½)
½�	½�	½�	½�	½*	½�½�½P   P   �	½Q	½�	½�	½.
½�	½�	½a
½Y
½-
½�	½U
½>
½7
½
½�	½'
½�	½�	½O	½P   P   O	½7	½=	½	½�	½
½�	½
½
½D
½�	½�	½:
½3
½
½�	½�	½�	½/	½O	½P   P   �	½�	½�	½,	½t	½n	½�	½t	½�	½ 
½/
½�	½L
½�	½�	½e	½�	½�	½F	½/	½P   P   �	½�	½�	½|	½�	½k	½�	½j	½�	½�	½�	½�	½�	½�	½�	½
½t	½�	½�	½�	½P   P   '
½�	½y	½�	½I
½
½�	½\	½�	½�	½j	½�	½�	½m	½�	½�	½k	½t	½�	½�	½P   P   �	½�	½(
½A
½�	½�	½�	½_	½�	½�	½�	½_	½�	½�	½`	½y	½�	½
½e	½�	½P   P   
½
½�
½;
½}
½8
½
½�	½�	½�	½�	½^	½	½_	½�½`	½�	½�	½�	½
½P   P   7
½}
½�
½�	½�	½�
½i
½B
½
½�	½�	½a	½�	½]	½_	½�	½m	½�	½�	½3
½P   P   >
½h
½�
½i
½�
½�
½�
½Y
½Q
½D
½<
½�	½�	½�	½	½�	½�	½�	½L
½:
½P   P   U
½�
½ ½�
½�½�½{
½ ½�
½B
½�	½�	½�	½a	½^	½_	½�	½�	½�	½�	½P   P   �	½S
½�
½�
½�
½0½½�
½�
½b
½�	½�	½<
½�	½�	½�	½j	½�	½/
½�	½P   P   -
½^
½½½�½�½�½�½½½b
½B
½D
½�	½�	½�	½�	½�	½ 
½D
½P   P   Y
½�
½�
½½?½4½/½$½Z½½�
½�
½Q
½
½�	½�	½�	½�	½�	½
½P   P   a
½=
½½�
½�½&½½O½$½�½�
½ ½Y
½B
½�	½_	½\	½j	½t	½
½P   P   �	½d
½�
½�
½�
½�½`½½/½�½½{
½�
½i
½
½�	½�	½�	½�	½�	½P   P   �	½@
½�
½k
½�½R½�½&½4½�½0½�½�
½�
½8
½�	½
½k	½n	½
½P   P   .
½�	½s
½�	½½�½�
½�½?½�½�
½�½�
½�	½}
½�	½I
½�	½t	½�	½P   P   �	½�	½3
½H
½�	½k
½�
½�
½½½�
½�
½i
½�	½;
½A
½�	½|	½,	½	½P   P   �	½�	½|	½3
½s
½�
½�
½½�
½½�
½ ½�
½�
½�
½(
½y	½�	½�	½=	½P   P   Q	½�	½�	½�	½�	½@
½d
½=
½�
½^
½S
½�
½h
½}
½
½�	½�	½�	½�	½7	½P   P   
½�	½�	½�	½�	½�	½�	½M
½j
½�
½�
½�
½\
½
½�	½	
½�	½�	½�	½�	½P   P   �	½�	½�	½
½
½�	½�
½7
½'
½K
½~
½O
½-
½[
½H
½�
½�	½$
½
½�	½P   P   �	½{	½�	½
½h
½�	½R
½W
½
½�	½�	½V
½
½�	½�	½W
½J
½�	½G
½
½P   P   �	½�	½�	½
½
½�	½�	½�	½1
½
½�	½k
½j
½�	½�	½>
½�	½�	½�	½$
½P   P   �	½
½U
½
½�	½�	½K
½�	½(
½�	½!
½�	½�	½�	½6
½�	½�	½�	½J
½�	½P   P   	
½�	½
½
½�	½
½�
½Y
½&
½�	½�	½

½�	½0
½%
½�	½�	½>
½W
½�
½P   P   �	½/
½
½)
½�	½Q
½�	½0
½
½
½&
½
½�
½�	½L
½%
½6
½�	½�	½H
½P   P   
½�
½z
½5½7½i
½�
½=
½F
½�	½�	½�	½
½h	½�	½0
½�	½�	½�	½[
½P   P   \
½�
½
½�	½�
½ 
½
½�
½Q
½H
½
½Q
½�	½
½�
½�	½�	½j
½
½-
½P   P   �
½�
½�
½3½�
½�
½½�
½�
½�
½]
½i
½Q
½�	½
½

½�	½k
½V
½O
½P   P   �
½�
½�
½T½�
½*
½½1½�
½�
½�
½]
½
½�	½&
½�	½!
½�	½�	½~
½P   P   �
½�
½�
½�
½�
½D½!½�
½�
½z
½�
½�
½H
½�	½
½�	½�	½
½�	½K
½P   P   j
½�
½�
½�
½t½½�½�
½^½�
½�
½�
½Q
½F
½
½&
½(
½1
½
½'
½P   P   M
½s
½�
½D½½�
½�
½�
½�
½�
½1½�
½�
½=
½0
½Y
½�	½�	½W
½7
½P   P   �	½�
½9
½%½�
½½�½�
½�½!½½½
½�
½�	½�
½K
½�	½R
½�
½P   P   �	½]
½q
½�	½�
½Q
½½�
½½D½*
½�
½ 
½i
½Q
½
½�	½�	½�	½�	½P   P   �	½�	½�	½.½½�
½�
½½t½�
½�
½�
½�
½7½�	½�	½�	½
½h
½
½P   P   �	½�	½

½I
½.½�	½%½D½�
½�
½T½3½�	½5½)
½
½
½
½
½
½P   P   �	½�	½�
½

½�	½q
½9
½�
½�
½�
½�
½�
½
½z
½
½
½U
½�	½�	½�	½P   P   �	½[	½�	½�	½�	½]
½�
½s
½�
½�
½�
½�
½�
½�
½/
½�	½
½�	½{	½�	½P   P   9	½
½ 
½2
½/
½�
½^
½|
½^
½!
½a
½=
½[
½S
½h
½�
½
½:
½
½
½P   P   
½"
½5
½�	½
½�	½
½!
½
½i
½�
½�
½W
½�
½>
½�	½�	½
½�	½K
½P   P   
½0
½

½�	½�	½`
½�	½�	½�
½�
½
½�	½
½�
½j
½�	½�	½]
½�	½�	½P   P   :
½?
½)
½E
½
½`
½�
½2
½�	½�	½A
½
½
½R
½
½�	½D
½�
½]
½
½P   P   
½
½�	½)
½
½�	½�	½B
½p
½�	½�
½E
½W
½1
½~
½
½Z
½D
½�	½�	½P   P   �
½ ½�
½}
½�
½�
½�	½�	½�	½
½\
½�	½�	½�	½�	½D
½
½�	½�	½�	½P   P   h
½v
½-
½1
½9
½
½H
½4
½j
½
½v
½�	½
½;
½�	½�	½~
½
½j
½>
½P   P   S
½u
½o
½�
½�
½f
½u
½z
½�
½�
½S
½9
½�	½
½;
½�	½1
½R
½�
½�
½P   P   [
½�
½�
½9½
½'½½�
½H
½k
½
½
½^
½�	½
½�	½W
½
½
½W
½P   P   =
½k
½-
½E½�
½�
½S½4
½o
½;
½~
½�	½
½9
½�	½�	½E
½
½�	½�
½P   P   a
½�
½�
½�
½,½�½½�
½½�
½U
½~
½
½S
½v
½\
½�
½A
½
½�
½P   P   !
½�
½7½�
½Y
½½½�
½½½�
½;
½k
½�
½
½
½�	½�	½�
½i
½P   P   ^
½}
½�
½½g½�½R½�½-½½½o
½H
½�
½j
½�	½p
½�	½�
½
½P   P   |
½�
½>
½�
½s
½o½/½>½�½�
½�
½4
½�
½z
½4
½�	½B
½2
½�	½!
½P   P   ^
½n
½½J½½½½/½R½½½S½½u
½H
½�	½�	½�
½�	½
½P   P   �
½y
½w
½,½�
½�½½o½�½½�½�
½'½f
½
½�
½�	½`
½`
½�	½P   P   /
½½1
½�
½)
½�
½½s
½g½Y
½,½�
½
½�
½9
½�
½
½
½�	½
½P   P   2
½
½t
½N
½�
½,½J½�
½½�
½�
½E½9½�
½1
½}
½)
½E
½�	½�	½P   P    
½0
½$
½t
½1
½w
½½>
½�
½7½�
½-
½�
½o
½-
½�
½�	½)
½

½5
½P   P   
½*
½0
½
½½y
½n
½�
½}
½�
½�
½k
½�
½u
½v
½ ½
½?
½0
½"
½P   P   H
½^
½�	½~
½Z
½
½�
½�
½�
½�
½g
½�
½�
½�
½�
½
½i
½�
½�	½[
½P   P   [
½i
½.
½d
½�
½�
½�
½}
½ 
½e
½�
½�
½v
½�	½�
½y
½�
½�
½Q
½F
½P   P   �	½f
½�	½a
½�	½U
½q
½�
½�
½W
½�
½�
½�
½Y
½v
½�
½�
½L
½
½Q
½P   P   �
½�
½�
½�
½�
½`
½�	½9
½�
½
½
½4
½8
½0
½6
½�
½/
½�	½L
½�
½P   P   i
½ 
½
½6
½O
½�
½b
½6
½J
½T
½$
½[
½�
½k
½�	½g
½]
½/
½�
½�
½P   P   
½�	½�
½}
½
½
½s
½�
½�
½
½_
½L
½�
½l
½b
½i
½g
½�
½�
½y
½P   P   �
½Q
½�
½�
½�
½=
½�
½�
½]
½9
½�	½\
½�
½F
½�
½b
½�	½6
½v
½�
½P   P   �
½C
½�
½V
½n
½�
½R
½�
½�	½w
½
½~
½�
½+
½F
½l
½k
½0
½Y
½�	½P   P   �
½�
½�
½½�
½�
½�
½�
½�
½u
½�
½J
½�
½�
½�
½�
½�
½8
½�
½v
½P   P   �
½(½�
½�	½�
½�
½
½�
½'½�
½�
½�
½J
½~
½\
½L
½[
½4
½�
½�
½P   P   g
½�
½½½�
½0½�
½
½&½�
½z
½�
½�
½
½�	½_
½$
½
½�
½�
½P   P   �
½�
½>
½�
½_½�
½�
½�½�
½/
½�
½�
½u
½w
½9
½
½T
½
½W
½e
½P   P   �
½½½�
½�
½�
½u
½�
½�
½�
½&½'½�
½�	½]
½�
½J
½�
½�
½ 
½P   P   �
½�
½�
½½]½�
½&½½�
½�½
½�
½�
½�
½�
½�
½6
½9
½�
½}
½P   P   �
½W
½�
½�	½�
½�
½]
½&½u
½�
½�
½
½�
½R
½�
½s
½b
½�	½q
½�
½P   P   
½5
½�
½½�
½½�
½�
½�
½�
½0½�
½�
½�
½=
½
½�
½`
½U
½�
½P   P   Z
½
½�
½P
½�
½�
½�
½]½�
½_½�
½�
½�
½n
½�
½
½O
½�
½�	½�
½P   P   ~
½.
½u
½�
½P
½½�	½½�
½�
½½�	½½V
½�
½}
½6
½�
½a
½d
½P   P   �	½�
½%
½u
½�
½�
½�
½�
½½>
½½�
½�
½�
½�
½�
½
½�
½�	½.
½P   P   ^
½s
½�
½.
½
½5
½W
½�
½½�
½�
½(½�
½C
½Q
½�	½ 
½�
½f
½i
½P   P   m
½_
½?
½2
½�
½r
½�
½�
½�
½�
½!½�
½�
½�
½�
½c
½�
½:
½:
½]
½P   P   ]
½h
½�
½�
½�	½p
½C
½�
½�
½�
½�	½&
½�
½�
½q
½G
½v
½�	½�
½�
½P   P   :
½M
½:
½�
½�
½f
½�
½`
½?
½e
½�
½�
½X
½s
½S
½q
½�
½Y
½�
½�
½P   P   :
½R
½S
½1
½�	½f
½�
½�
½v
½�
½�
½U
½X
½�
½�
½c
½�
½�
½Y
½�	½P   P   �
½�
½�
½�
½�
½{
½�
½�
½�	½p
½x
½T
½
½�
½k
½w
½
½�
½�
½v
½P   P   c
½T
½d
½Q
½�
½o
½$
½x
½b
½�
½M
½�
½I
½
½�
½f
½w
½c
½q
½G
½P   P   �
½(½�
½d
½�
½�
½�
½�
½=
½�
½g
½�
½=
½
½�
½�
½k
½�
½S
½q
½P   P   �
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½<
½1
½
½
½�
½�
½s
½�
½P   P   �
½>
½�
½�
½_½[
½�
½A
½�
½�
½W
½|
½�	½<
½=
½I
½
½X
½X
½�
½P   P   �
½
½R½½�
½½=½C½
½�
½
½�
½|
½�
½�
½�
½T
½U
½�
½&
½P   P   !½½d
½�
½�
½w
½�
½�
½p
½�
½<½
½W
½�
½g
½M
½x
½�
½�
½�	½P   P   �
½�
½½�
½@½$½,½G½�
½ ½�
½�
½�
½�
½�
½�
½p
½�
½e
½�
½P   P   �
½�	½�
½�
½�
½�
½�½�
½�
½�
½p
½
½�
½�
½=
½b
½�	½v
½?
½�
½P   P   �
½^
½i½�
½,½½5½½�
½G½�
½C½A
½�
½�
½x
½�
½�
½`
½�
½P   P   �
½�
½�
½½½>½V½5½�½,½�
½=½�
½�
½�
½$
½�
½�
½�
½C
½P   P   r
½½�
½�
½½1
½>½½�
½$½w
½½[
½�
½�
½o
½{
½f
½f
½p
½P   P   �
½~
½�
½�
½3½½½,½�
½@½�
½�
½_½�
½�
½�
½�
½�	½�
½�	½P   P   2
½�
½K
½�
½�
½�
½½�
½�
½�
½�
½½�
½�
½d
½Q
½�
½1
½�
½�
½P   P   ?
½H
½�
½K
½�
½�
½�
½i½�
½½d
½R½�
½�
½�
½d
½�
½S
½:
½�
½P   P   _
½W
½H
½�
½~
½½�
½^
½�	½�
½½
½>
½�
½(½T
½�
½R
½M
½h
½P   P   ]
½n
½+½�
½�
½�
½H
½z
½�
½�
½{
½�
½�
½�
½F
½�
½�
½�
½-½o
½P   P   o
½�
½
½"
½Q
½�
½�
½�
½½�
½�
½�
½�
½�
½�
½�
½�
½4
½,
½
½P   P   -½�
½½<
½�
½�
½U
½
½y
½�
½�
½�
½w
½�
½�
½�
½>
½�
½�
½,
½P   P   �
½M
½k
½�
½H
½�
½�
½�
½n
½�
½�
½�
½�
½�
½�
½b
½�
½�
½�
½4
½P   P   �
½~
½z
½n
½�
½�
½`
½�
½�
½�
½E
½�
½�
½�
½Y
½�
½�
½�
½>
½�
½P   P   �
½�
½�
½�
½�
½�
½�
½z
½`
½�
½�
½�
½�
½�
½[
½�
½�
½b
½�
½�
½P   P   F
½�
½�
½�
½s
½b
½e
½�
½�
½�
½X
½`
½(
½½~
½[
½Y
½�
½�
½�
½P   P   �
½�
½�
½�
½½�
½�
½�
½�
½�
½~
½�
½�
½F½½�
½�
½�
½�
½�
½P   P   �
½�
½�
½g
½p
½I
½�
½�
½�
½�
½�
½�
½�
½�
½(
½�
½�
½�
½w
½�
½P   P   �
½�
½�
½½�
½�
½½�
½½�
½�
½�
½�
½�
½`
½�
½�
½�
½�
½�
½P   P   {
½�
½�
½
½½½½
½�
½�
½�
½�
½�
½~
½X
½�
½E
½�
½�
½�
½P   P   �
½m
½Y½½e
½�
½�
½a
½ ½l½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½P   P   �
½�
½�
½
½_½�
½�
½�
½^½ ½�
½½�
½�
½�
½`
½�
½n
½y
½½P   P   z
½½�
½�	½X
½�
½�
½�
½�
½a
½
½�
½�
½�
½�
½z
½�
½�
½
½�
½P   P   H
½�
½�
½�
½:½�
½�
½�
½�
½�
½½½�
½�
½e
½�
½`
½�
½U
½�
½P   P   �
½�
½�
½�
½�
½�
½�
½�
½�
½�
½½�
½I
½�
½b
½�
½�
½�
½�
½�
½P   P   �
½�
½b
½ ½+
½�
½:½X
½_½e
½½�
½p
½½s
½�
½�
½H
½�
½Q
½P   P   �
½|
½�
½�
½ ½�
½�
½�	½
½½
½½g
½�
½�
½�
½n
½�
½<
½"
½P   P   +½X
½w
½�
½b
½�
½�
½�
½�
½Y½�
½�
½�
½�
½�
½�
½z
½k
½½
½P   P   n
½�
½X
½|
½�
½�
½�
½½�
½m
½�
½�
½�
½�
½�
½�
½~
½M
½�
½�
½P   P   4½�
½�
½�
½t
½n
½�
½�
½V
½�
½�
½�
½r
½�
½�
½o
½Y
½�
½�
½�
½P   P   �
½�
½�
½�
½½�
½�
½�
½9
½�
½�
½�
½x
½$
½�
½�
½�
½½�
½�
½P   P   �
½�	½�
½�
½�
½�
½�
½�
½�
½�
½�
½w
½�
½�
½�
½�
½�
½{
½�
½�
½P   P   �
½�
½�
½�
½½o
½f
½
½�
½�
½�
½�
½t
½�
½�
½�
½�
½w
½{
½½P   P   Y
½B
½�
½#
½U
½�
½�
½�
½�
½�
½l
½i
½n
½�
½v
½�
½�
½�
½�
½�
½P   P   o
½�
½�
½�
½�
½t
½�
½�
½�
½�
½�
½�
½�
½q
½�
½�
½�
½�
½�
½�
½P   P   �
½�
½�
½�
½�
½t
½�
½�
½�
½�
½x
½�
½V
½"
½o
½�
½v
½�
½�
½�
½P   P   �
½�
½ ½�
½�
½�
½½�
½
½�
½�
½}
½v
½9
½"
½q
½�
½�
½�
½$
½P   P   r
½�
½x
½i½�
½n½|
½�
½
½�
½�
½�
½g
½v
½V
½�
½n
½t
½�
½x
½P   P   �
½:½@
½�
½�
½�
½�
½N
½M½�
½�
½U
½�
½}
½�
½�
½i
½�
½w
½�
½P   P   �
½�
½\½t½2½�
½1½o½I½�
½�
½�
½�
½�
½x
½�
½l
½�
½�
½�
½P   P   �
½�
½�	½�
½!½�
½�
½/½�
½�	½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½P   P   V
½3½N½�
½½�
½�
½�
½�
½�
½I½M½
½
½�
½�
½�
½�
½�
½9
½P   P   �
½�
½U
½n½-½�
½R½Z½�
½/½o½N
½�
½�
½�
½�
½�
½
½�
½�
½P   P   �
½½U
½�
½5½�
½½R½�
½�
½1½�
½|
½½�
½�
½�
½f
½�
½�
½P   P   n
½�
½�
½�½�
½�
½�
½�
½�
½�
½�
½�
½n½�
½t
½t
½�
½o
½�
½�
½P   P   t
½�
½�
½�
½�
½�
½5½-½½!½2½�
½�
½�
½�
½�
½U
½½�
½½P   P   �
½$
½�
½�
½�
½�½�
½n½�
½�
½t½�
½i½�
½�
½�
½#
½�
½�
½�
½P   P   �
½�
½�
½�
½�
½�
½U
½U
½N½�	½\½@
½x
½ ½�
½�
½�
½�
½�
½�
½P   P   �
½�	½�
½$
½�
½�
½½�
½3½�
½�
½:½�
½�
½�
½�
½B
½�
½�	½�
½P   P   
½�
½7
½j
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½Z
½V
½�
½P   P   �
½�
½½�
½�
½x
½q
½p
½6½*½�
½t
½½M½�
½W
½�
½�
½�
½½P   P   V
½�
½A
½�
½a
½�
½�
½:
½�
½�
½�
½�
½�
½�
½�
½4
½½�
½E
½�
½P   P   Z
½�
½½b
½�
½�
½3½�
½�
½�
½�
½½½�
½�
½�
½�
½+½�
½�
½P   P   �
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½
½�
½½�
½P   P   �
½P½M
½V
½E½�
½r
½8
½�
½�
½}
½g
½�
½�
½}
½m
½�
½�
½4
½W
½P   P   �
½�
½�
½�
½�
½�
½�
½
½�
½�
½�
½x
½½	½�
½}
½�
½�
½�
½�
½P   P   �
½�
½N
½k
½F
½H
½�
½�
½<½�
½�
½�
½�
½�
½	½�
½�
½�
½�
½M½P   P   �
½�
½½�
½�
½½
½�
½½!½�
½½�
½�
½½�
½�
½½�
½½P   P   �
½%
½�
½�
½�
½�
½�
½�
½*
½�
½j
½�
½½�
½x
½g
½�
½½�
½t
½P   P   �
½ ½�
½½E
½�
½>
½½�
½ ½½j
½�
½�
½�
½}
½�
½�
½�
½�
½P   P   �
½@½½�
½�
½½½�
½�
½�
½ ½�
½!½�
½�
½�
½�
½�
½�
½*½P   P   �
½6
½�
½�
½�
½�
½�
½�
½}
½�
½�
½*
½½<½�
½�
½�
½�
½�
½6½P   P   �
½�
½�
½)½�
½�
½�
½�
½�
½�
½½�
½�
½�
½
½8
½�
½�
½:
½p
½P   P   �
½�
½½�
½
½�
½�
½�
½�
½½>
½�
½
½�
½�
½r
½�
½3½�
½q
½P   P   �
½�
½B
½�
½�
½*½�
½�
½�
½½�
½�
½½H
½�
½�
½�
½�
½�
½x
½P   P   �
½7½�
½X
½�
½�
½
½�
½�
½�
½E
½�
½�
½F
½�
½E½�
½�
½a
½�
½P   P   j
½�
½\
½�
½X
½�
½�
½)½�
½�
½½�
½�
½k
½�
½V
½�
½b
½�
½�
½P   P   7
½½�
½\
½�
½B
½½�
½�
½½�
½�
½½N
½�
½M
½�
½½A
½½P   P   �
½�
½½�
½7½�
½�
½�
½6
½@½ ½%
½�
½�
½�
½P½�
½�
½�
½�
½P   P   8
½�
½�
½�
½�
½�
½�
½P
½�
½�
½�
½ ½�
½2
½�
½�
½�
½�
½�
½�
½P   P   �
½�
½w
½�
½�
½�
½�
½�
½�
½x
½.½�
½f
½�
½�
½�
½�
½�
½�
½v
½P   P   �
½?½�
½�
½�
½�
½�
½�
½�
½S
½�
½�
½�
½]
½�
½�
½�
½�
½�
½�
½P   P   �
½X
½M
½�
½�
½�
½.
½�
½�
½d
½e
½z
½�
½Z
½h
½½�
½,
½�
½�
½P   P   �
½½y
½�
½�
½�
½�
½�
½½�
½½�
½�
½�
½½�
½�
½�
½�
½�
½P   P   �
½$
½�
½�
½
½�
½½�
½�
½�
½�
½u
½�
½�
½�
½�
½�
½½�
½�
½P   P   �
½�
½�
½s½�
½�
½�
½�
½�
½�
½�
½�
½�
½F
½�
½�
½½h
½�
½�
½P   P   2
½�
½�
½P½?½�
½�
½B
½�
½9
½p
½�
½�
½)
½F
½�
½�
½Z
½]
½�
½P   P   �
½�
½�
½U
½�
½m
½�
½�
½�
½
½�
½w
½�
½�
½�
½�
½�
½�
½�
½f
½P   P    ½½8½�
½½�
½�
½`½ ½�
½½½w
½�
½�
½u
½�
½z
½�
½�
½P   P   �
½v
½l
½�
½�
½+½�
½�
½X
½�
½�
½½�
½p
½�
½�
½½e
½�
½.½P   P   �
½�
½s½½�
½�
½�
½�
½½j½�
½�
½
½9
½�
½�
½�
½d
½S
½x
½P   P   �
½(½M
½�
½½2½�
½(½½½X
½ ½�
½�
½�
½�
½½�
½�
½�
½P   P   P
½�
½*½�
½½½�
½
½(½�
½�
½`½�
½B
½�
½�
½�
½�
½�
½�
½P   P   �
½�
½½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½½�
½.
½�
½�
½P   P   �
½�
½�
½3
½�
½j½�
½½2½�
½+½�
½m
½�
½�
½�
½�
½�
½�
½�
½P   P   �
½
½�
½K½�
½�
½�
½½½�
½�
½½�
½?½�
½
½�
½�
½�
½�
½P   P   �
½�
½�
½V½K½3
½�
½�
½�
½½�
½�
½U
½P½s½�
½�
½�
½�
½�
½P   P   �
½L
½�
½�
½�
½�
½½*½M
½s½l
½8½�
½�
½�
½�
½y
½M
½�
½w
½P   P   �
½W½L
½�
½
½�
½�
½�
½(½�
½v
½½�
½�
½�
½$
½½X
½?½�
½P   P   �½�
½�
½�
½�
½�
½�
½/½�
½�
½�
½�
½�
½(½�
½�
½�
½�
½�
½�
½P   P   �
½s
½r
½�
½I
½�
½l
½�
½�
½y
½�
½�
½
½�
½�
½�
½�
½@
½�
½v
½P   P   �
½R
½½�
½�
½�
½�
½�
½�
½x½½K
½&½q½�
½�
½~
½�
½�
½�
½P   P   �
½�
½�
½�
½\
½�
½�
½�
½e
½�
½	½�
½�
½�
½�
½y
½�
½�
½�
½@
½P   P   �
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½
½�
½~
½�
½P   P   �
½�
½-½=½�
½�
½�
½�
½t
½x
½�
½�
½�
½�
½�
½�
½�
½y
½�
½�
½P   P   �
½�
½|
½�	½i
½�
½�
½�
½�
½�
½�
½�
½½�
½½�
½�
½�
½�
½�
½P   P   (½.½N½\
½c
½W½½6½�
½_½½�
½�
½�
½�
½�
½�
½�
½q½�
½P   P   �
½a
½=
½�
½�
½�
½F
½v
½�
½�
½½�
½½�
½½�
½�
½�
½&½
½P   P   �
½'½�
½�
½�
½�
½�
½�
½½
½�
½b
½�
½�
½�
½�
½�
½�
½K
½�
½P   P   �
½�
½�
½�
½"½
½<½�
½�
½�
½�
½�
½½½�
½�
½�
½	½½�
½P   P   �
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½
½�
½_½�
½x
½�
½�
½x½y
½P   P   �
½@½�
½|
½A
½�
½�
½�
½Z
½�
½�
½½�
½�
½�
½t
½�
½e
½�
½�
½P   P   /½D
½b
½�
½�
½�
½½½�
½�
½�
½�
½v
½6½�
½�
½�
½�
½�
½�
½P   P   �
½½z
½�
½ ½�
½�
½½�
½�
½<½�
½F
½½�
½�
½�
½�
½�
½l
½P   P   �
½�
½V½�
½�
½,
½�
½�
½�
½�
½
½�
½�
½W½�
½�
½�
½�
½�
½�
½P   P   �
½�
½r
½d
½½�
½ ½�
½A
½�
½"½�
½�
½c
½i
½�
½�
½\
½�
½I
½P   P   �
½�
½3½�	½d
½�
½�
½�
½|
½�
½�
½�
½�
½\
½�	½=½�
½�
½�
½�
½P   P   �
½�
½�
½3½r
½V½z
½b
½�
½�
½�
½�
½=
½N½|
½-½�
½�
½½r
½P   P   �
½Y
½�
½�
½�
½�
½½D
½@½�
½�
½'½a
½.½�
½�
½�
½�
½R
½s
½P   P   �
½�
½�
½{
½�
½ ½:
½½�
½�
½#½�
½�
½0½*
½�
½�
½�
½�
½�
½P   P   �
½�
½
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½½P   P   �
½�
½�
½�
½�
½�
½�
½�
½[
½s
½}
½�
½�
½_
½�
½�
½�
½�
½�
½�
½P   P   �
½!½½�
½ ½�
½�
½�
½�
½�
½%
½�
½�
½
½�
½�
½�
½½�
½�
½P   P   �
½�	½I
½
½�
½�
½�
½�
½�
½@½m
½�
½�
½�
½�
½&½�
½�
½�
½�
½P   P   �
½½�
½
½�
½�
½�
½�
½�
½½�
½�
½t
½�
½�
½�
½&½�
½�
½�
½P   P   *
½C
½½.½½P
½,
½�
½j
½�
½�
½�
½^
½�
½h
½�
½�
½�
½�
½�
½P   P   0½�
½?
½�
½�
½=
½a
½.½�
½l
½3
½�
½r
½�
½�
½�
½�
½
½_
½�
½P   P   �
½�
½�
½�
½�
½�
½½�
½�
½�
½�
½�
½�
½r
½^
½t
½�
½�
½�
½�
½P   P   �
½N
½�
½�
½�
½�
½�
½�
½N
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½�
½P   P   #½�
½
½k
½�
½�
½{
½�
½ ½�
½�
½�
½�
½3
½�
½�
½m
½%
½}
½�
½P   P   �
½�
½�
½½�
½½½�
½�
½�
½�
½�
½�
½l
½�
½½@½�
½s
½�
½P   P   �
½d
½"½
½=½�
½(½�
½M½�
½ ½N
½�
½�
½j
½�
½�
½�
½[
½�
½P   P   ½�
½�
½s
½�
½�
½
½j
½�
½�
½�
½�
½�
½.½�
½�
½�
½�
½�
½�
½P   P   :
½r
½½�
½�
½$½½
½(½½{
½�
½½a
½,
½�
½�
½�
½�
½�
½P   P    ½>
½M
½�
½�
½�
½$½�
½�
½½�
½�
½�
½=
½P
½�
½�
½�
½�
½�
½P   P   �
½½½�
½�
½�
½�
½�
½=½�
½�
½�
½�
½�
½½�
½�
½ ½�
½�
½P   P   {
½ 
½�
½3½�
½�
½�
½s
½
½½k
½�
½�
½�
½.½
½
½�
½�
½�
½P   P   �
½%½"
½�
½½M
½½�
½"½�
½
½�
½�
½?
½½�
½I
½½�
½
½P   P   �
½�
½%½ 
½½>
½r
½�
½d
½�
½�
½N
½�
½�
½C
½½�	½!½�
½�
½P   P   �	½�
½"
½�
½u
½u
½½
½�
½�
½�
½x
½�
½B
½½\
½�
½�
½
½�
½P   P   �
½�
½�
½�
½!½l
½�
½�
½�
½�
½�
½�
½½Y
½�
½�
½T
½½�
½�
½P   P   
½�
½,
½�
½�
½8
½o
½�
½�
½�
½�
½½�
½}
½½�
½w
½O
½z
½�
½P   P   �
½�
½�
½�
½½Q
½�
½k
½�
½�
½�
½�
½�
½�
½�
½d
½]
½�
½O
½½P   P   �
½"½-½0½�
½I
½}
½H
½k
½u
½�
½�
½	
½�
½�
½T
½�
½]
½w
½T
½P   P   \
½�
½s
½k
½f
½`
½�
½�
½�
½N
½\
½½�
½
½�
½�
½T
½d
½�
½�
½P   P   ½½�
½�
½�
½½½�
½�
½�
½�
½�
½]
½�
½f
½�
½�
½�
½½�
½P   P   B
½�
½�
½�
½�
½�
½�
½$
½�
½�
½�
½�
½�
½�
½�
½
½�
½�
½}
½Y
½P   P   �
½�
½�
½k
½G
½d
½�
½�
½�
½�
½�
½�
½4
½�
½]
½�
½	
½�
½�
½½P   P   x
½�
½�
½j
½�
½�
½�
½�
½�
½�
½�
½½�
½�
½�
½½�
½�
½½�
½P   P   �
½�
½�
½�
½�
½½�
½�
½�
½�
½
½�
½�
½�
½�
½\
½�
½�
½�
½�
½P   P   �
½�
½&
½�
½�
½*
½K
½�
½t
½;
½�
½�
½�
½�
½�
½N
½u
½�
½�
½�
½P   P   �
½�
½�
½�
½�
½x
½�
½�
½�
½t
½�
½�
½�
½�
½�
½�
½k
½�
½�
½�
½P   P   
½�
½�
½�
½
½�
½�
½�
½�
½�
½�
½�
½�
½$
½�
½�
½H
½k
½�
½�
½P   P   ½�
½�
½}
½�
½U
½p
½�
½�
½K
½�
½�
½�
½�
½½�
½}
½�
½o
½�
½P   P   u
½�
½�
½s
½�
½�
½U
½�
½x
½*
½½�
½d
½�
½½`
½I
½Q
½8
½l
½P   P   u
½i
½�
½�
½A
½�
½�
½
½�
½�
½�
½�
½G
½�
½�
½f
½�
½½�
½!½P   P   �
½I½y
½�
½�
½s
½}
½�
½�
½�
½�
½j
½k
½�
½�
½k
½0½�
½�
½�
½P   P   "
½�
½�
½y
½�
½�
½�
½�
½�
½&
½�
½�
½�
½�
½�
½s
½-½�
½,
½�
½P   P   �
½�
½�
½I½i
½�
½�
½�
½�
½�
½�
½�
½�
½�
½½�
½"½�
½�
½�
½P   P   �
½�
½�
½�
½h
½x
½�
½�
½�
½�
½�
½X
½�
½�
½�
½s
½t
½�
½�
½�
½P   P   �
½�
½_
½�
½W
½�
½>
½{
½�
½n
½{
½�
½�
½�
½k
½<
½�
½T
½�
½d
½P   P   �
½½�
½�
½Y
½�
½�
½+
½�
½�
½n
½I
½R
½�
½�
½&
½�
½�
½H
½�
½P   P   �
½
½
½�
½D
½�
½½�
½z
½W
½�
½�
½�
½�
½j
½a
½�
½�
½�
½T
½P   P   t
½�
½B
½�
½�
½�
½�
½�
½F½�
½L
½@
½�
½I
½
½�
½l½�
½�
½�
½P   P   s
½�
½�
½�
½v
½\
½K
½%
½�
½|
½�
½J
½�
½�
½D
½½�
½a
½&
½<
½P   P   �
½�
½]
½X
½[
½�
½�
½�
½�
½E
½`
½N
½W
½�
½U
½D
½
½j
½�
½k
½P   P   �
½[
½�
½�
½�
½�
½k
½|
½�
½�
½�
½,
½�
½�
½�
½�
½I
½�
½�
½�
½P   P   �
½y
½X
½½ ½½;
½�
½�
½c
½f
½�
½�
½�
½W
½�
½�
½�
½R
½�
½P   P   X
½�
½X
½x
½�
½y
½�
½E
½�
½w
½�
½N
½�
½,
½N
½J
½@
½�
½I
½�
½P   P   �
½�
½�
½�
½�
½
½�
½�
½�
½�
½�
½�
½f
½�
½`
½�
½L
½�
½n
½{
½P   P   �
½�
½�
½�
½½�
½�
½�
½�
½�
½�
½w
½c
½�
½E
½|
½�
½W
½�
½n
½P   P   �
½�
½�
½�
½4
½�
½�
½�
½c
½�
½�
½�
½�
½�
½�
½�
½F½z
½�
½�
½P   P   �
½�
½J
½�
½�
½�
½�
½m
½�
½�
½�
½E
½�
½|
½�
½%
½�
½�
½+
½{
½P   P   �
½p
½3
½�
½�
½�
½�
½�
½�
½�
½�
½�
½;
½k
½�
½K
½�
½½�
½>
½P   P   x
½�
½�
½½�
½
½�
½�
½�
½�
½
½y
½½�
½�
½\
½�
½�
½�
½�
½P   P   h
½t
½g
½�
½�
½�
½�
½�
½4
½½�
½�
½ ½�
½[
½v
½�
½D
½Y
½W
½P   P   �
½�
½�
½D
½�
½½�
½�
½�
½�
½�
½x
½½�
½X
½�
½�
½�
½�
½�
½P   P   �
½
½,
½�
½g
½�
½3
½J
½�
½�
½�
½X
½X
½�
½]
½�
½B
½
½�
½_
½P   P   �
½½
½�
½t
½�
½p
½�
½�
½�
½�
½�
½y
½[
½�
½�
½�
½
½½�
½P   P   �½
½�
½m
½�
½�
½D
½�
½1
½q
½}
½Z
½ 
½�
½U
½�
½�
½g
½�
½
½P   P   
½
½
½�
½
½�
½s
½�
½\
½}
½�
½	½�
½s
½�
½]
½�
½
½�
½
½P   P   �
½F
½�
½�
½�
½T
½W
½�
½
½d
½�
½l
½n
½N
½q
½�
½g
½_
½�
½�
½P   P   g
½�
½�
½l
½
½T
½�	½B
½�
½�
½d
½�
½�
½�
½�
½�
½I
½u	½_
½
½P   P   �
½5
½<
½%
½�
½�
½W
½@
½
½�
½�
½}
½½x
½}
½�
½�	½I
½g
½�
½P   P   �
½�
½�
½�
½�
½�
½g
½�
½�
½�
½�
½�
½^
½e
½�
½�
½�
½�
½�
½]
½P   P   U
½
½�
½ ½�
½/
½P
½�
½z
½�
½�
½�
½�
½O
½�
½�
½}
½�
½q
½�
½P   P   �
½N
½w
½V
½V
½e
½W
½�
½c
½\
½r
½o
½d
½>
½O
½e
½x
½�
½N
½s
½P   P    
½�
½�
½Q
½Z
½~
½�
½�
½5
½�
½�
½�
½½d
½�
½^
½½�
½n
½�
½P   P   Z
½v
½�
½�
½�
½X
½�
½�
½g
½b
½�
½j
½�
½o
½�
½�
½}
½�
½l
½	½P   P   }
½P
½'
½7
½%
½�
½[
½9
½*
½@
½�
½�
½�
½r
½�
½�
½�
½d
½�
½�
½P   P   q
½J
½w
½�
½
½�
½�
½�	½�
½�
½@
½b
½�
½\
½�
½�
½�
½�
½d
½}
½P   P   1
½_
½6
½�
½�
½�
½p
½�
½�
½�
½*
½g
½5
½c
½z
½�
½
½�
½
½\
½P   P   �
½�
½�
½1
½
½�
½C
½Z
½�
½�	½9
½�
½�
½�
½�
½�
½@
½B
½�
½�
½P   P   D
½L
½�
½�
½3
½�
½m
½C
½p
½�
½[
½�
½�
½W
½P
½g
½W
½�	½W
½s
½P   P   �
½9
½a
½h
½|
½�
½�
½�
½�
½�
½�
½X
½~
½e
½/
½�
½�
½T
½T
½�
½P   P   �
½�
½�
½g
½D
½|
½3
½
½�
½
½%
½�
½Z
½V
½�
½�
½�
½
½�
½
½P   P   m
½%
½�
½½g
½h
½�
½1
½�
½�
½7
½�
½Q
½V
½ ½�
½%
½l
½�
½�
½P   P   �
½�
½A
½�
½�
½a
½�
½�
½6
½w
½'
½�
½�
½w
½�
½�
½<
½�
½�
½
½P   P   
½:
½�
½%
½�
½9
½L
½�
½_
½J
½P
½v
½�
½N
½
½�
½5
½�
½F
½
½P   P   L
½�
½q
½a
½�
½>
½z
½V
½W
½�
½
½�
½3
½#
½�
½i
½�
½X
½t
½�
½P   P   �
½�
½�
½�	½�
½�	½b
½,
½F
½�
½�	½�	½�
½{
½>
½B
½�	½�
½�	½�
½P   P   t
½�	½V
½
½�
½�
½�
½_
½
½�
½s
½u
½y
½�
½�	½j
½�
½�
½�
½�	½P   P   X
½L
½\
½l
½�
½�
½½�
½l
½�
½<
½
½
½C
½�
½z
½�
½½�
½�
½P   P   �
½h
½½\
½�
½�	½�
½�
½1
½A
½�
½�
½�	½�
½}
½\
½
½�
½�
½�	½P   P   i
½P
½"
½"
½N
½^
½E
½o
½H
½^
½�	½1
½:
½F
½J
½r	½\
½z
½j
½B
½P   P   �
½l
½T
½�	½^
½�
½}
½*
½
½�
½g
½=
½�
½j
½�
½J
½}
½�
½�	½>
½P   P   #
½�
½�
½n
½h
½�
½�
½K
½X
½�
½J
½�
½H
½I
½j
½F
½�
½C
½�
½{
½P   P   3
½
½1
½
½�
½/
½O
½�	½D
½�
½y
½
½�	½H
½�
½:
½�	½
½y
½�
½P   P   �
½�
½G
½�
½�
½|
½V
½e
½�
½�
½�	½n
½
½�
½=
½1
½�
½
½u
½�	½P   P   
½�
½p
½�
½[
½�
½�
½�
½}
½�
½
½�	½y
½J
½g
½�	½�
½<
½s
½�	½P   P   �
½�
½R
½~
½t
½u
½N
½r
½y
½A
½�
½�
½�
½�
½�
½^
½A
½�
½�
½�
½P   P   W
½�
½~
½q
½�
½t
½�	½_
½�
½y
½}
½�
½D
½X
½
½H
½1
½l
½
½F
½P   P   V
½�	½e
½�
½�
½]
½�
½*½_
½r
½�
½e
½�	½K
½*
½o
½�
½�
½_
½,
½P   P   z
½�
½Z
½a
½�
½=
½
½�
½�	½N
½�
½V
½O
½�
½}
½E
½�
½½�
½b
½P   P   >
½�
½�
½
½�
½�
½=
½]
½t
½u
½�
½|
½/
½�
½�
½^
½�	½�
½�
½�	½P   P   �
½V
½=
½p
½�
½�
½�
½�
½�
½t
½[
½�
½�
½h
½^
½N
½�
½�
½�
½�
½P   P   a
½D
½(
½�	½p
½
½a
½�
½q
½~
½�
½�
½
½n
½�	½"
½\
½l
½
½�	½P   P   q
½W
½½(
½=
½�
½Z
½e
½~
½R
½p
½G
½1
½�
½T
½"
½½\
½V
½�
½P   P   �
½�	½W
½D
½V
½�
½�
½�	½�
½�
½�
½�
½
½�
½l
½P
½h
½L
½�	½�
½P   P   �½H
½U
½\
½L
½
½3
½N
½�
½%
½�
½G
½�
½
½?
½4
½
½W
½Z
½G
½P   P   G
½P
½'
½9
½�
½8
½�
½O
½z
½�	½b
½I
½�	½�
½h
½�
½H
½�
½7
½'
½P   P   Z
½�
½N
½;
½�	½�	½>
½�	½�
½C
½9
½�
½L
½F
½m
½�	½>
½�	½�	½7
½P   P   W
½�	½�	½[
½�
½�	½$
½�	½a
½�	½
½r
½x
½�	½�	½e
½�	½)
½�	½�
½P   P   
½'
½'
½.
½)
½S
½4
½�	½�
½�
½[
½�
½O
½�
½c
½�
½�
½�	½>
½H
½P   P   4
½�
½�
½�
½k
½.
½�
½�	½0
½�
½�
½>
½b
½i
½Y
½�
½�
½e
½�	½�
½P   P   ?
½�	½J
½?
½j
½

½:
½O
½�
½
½4
½J
½�	½`
½�	½Y
½c
½�	½m
½h
½P   P   
½:
½)
½�
½{
½
½2
½C
½�
½,
½
½�
½n
½?
½`
½i
½�
½�	½F
½�
½P   P   �
½�
½E
½\
½f
½b
½c
½l
½�
½�	½=
½w
½5
½n
½�	½b
½O
½x
½L
½�	½P   P   G
½9
½�	½l
½#
½,
½Y
½�	½:
½+
½Z
½�
½w
½�
½J
½>
½�
½r
½�
½I
½P   P   �
½�	½F
½Z
½ 
½�	½
½3
½K
½
½�
½Z
½=
½
½4
½�
½[
½
½9
½b
½P   P   %
½�	½V
½
½Y
½�
½�
½�
½%
½,
½
½+
½�	½,
½
½�
½�
½�	½C
½�	½P   P   �
½A
½=
½
½ 
½d
½$
½P
½�	½%
½K
½:
½�
½�
½�
½0
½�
½a
½�
½z
½P   P   N
½a
½
½6
½�
½+
½�	½+
½P
½�
½3
½�	½l
½C
½O
½�	½�	½�	½�	½O
½P   P   3
½(
½`
½U
½"
½�
½{
½�	½$
½�
½
½Y
½c
½2
½:
½�
½4
½$
½>
½�
½P   P   
½
½"
½^
½
½�	½�
½+
½d
½�
½�	½,
½b
½
½

½.
½S
½�	½�	½8
½P   P   L
½{
½K
½p
½�
½
½"
½�
½ 
½Y
½ 
½#
½f
½{
½j
½k
½)
½�
½�	½�
½P   P   \
½
½�
½^
½p
½^
½U
½6
½
½
½Z
½l
½\
½�
½?
½�
½.
½[
½;
½9
½P   P   U
½�	½C
½�
½K
½"
½`
½
½=
½V
½F
½�	½E
½)
½J
½�
½'
½�	½N
½'
½P   P   H
½�
½�	½
½{
½
½(
½a
½A
½�	½�	½9
½�
½:
½�	½�
½'
½�	½�
½P
½P   P   �½%
½�	½)
½�	½
½
½�	½
½
½�
½
½"
½�	½
½
½�	½0
½�	½"
½P   P   "
½
½�	½�
½�	½>
½
½�	½�	½
½X
½Y
½
½�	½	
½
½P
½�	½�
½�	½P   P   �	½
½�	½�
½
½i
½E
½(
½h
½*
½B
½F	½C
½@
½Z
½0
½N
½Z
½$
½�
½P   P   0
½�
½{
½
½�	½d
½?
½L
½w
½
½�
½�	½�	½}
½
½p
½M
½?
½Z
½�	½P   P   �	½/
½�	½I
½�	½P
½8
½W
½
½[	½

½�	½)
½�	½

½p	½
½M
½N
½P
½P   P   
½L
½
½�	½C
½
½
½C
½X
½|	½p
½
½"
½
½
½X
½p	½p
½0
½
½P   P   
½P
½	
½'
½	
½E
½
½�	½[
½
½�	½
½)
½+
½*
½
½

½
½Z
½	
½P   P   �	½
½�	½ 
½	
½
½!
½�	½�	½7
½
½�	½#
½
½+
½
½�	½}
½@
½�	½P   P   "
½h
½H
½ 
½n	½�	½?
½T
½,
½
½5
½�	½
½#
½)
½"
½)
½�	½C
½
½P   P   
½
½.
½F
½i
½�
½c
½A
½
½�	½]
½G	½�	½�	½
½
½�	½�	½F	½Y
½P   P   �
½�	½�
½�	½0
½�
½�	½�	½w
½�	½�
½]
½5
½
½�	½p
½

½�
½B
½X
½P   P   
½�	½�
½+
½�	½
½
½(
½P
½y
½�	½�	½
½7
½
½|	½[	½
½*
½
½P   P   
½
½n
½<
½�
½0
½;
½'
½*
½P
½w
½
½,
½�	½[
½X
½
½w
½h
½�	½P   P   �	½U
½I
½�	½ 
½�	½3
½5
½'
½(
½�	½A
½T
½�	½�	½C
½W
½L
½(
½�	½P   P   
½'
½9
½J
½'
½
½e
½3
½;
½
½�	½c
½?
½!
½
½
½8
½?
½E
½
½P   P   
½C
½�	½
½x
½~
½
½�	½0
½
½�
½�
½�	½
½E
½
½P
½d
½i
½>
½P   P   �	½Q
½
½�	½�	½x
½'
½ 
½�
½�	½0
½i
½n	½	
½	
½C
½�	½�	½
½�	½P   P   )
½2
½�	½I
½�	½
½J
½�	½<
½+
½�	½F
½ 
½ 
½'
½�	½I
½
½�
½�
½P   P   �	½{
½�	½�	½
½�	½9
½I
½n
½�
½�
½.
½H
½�	½	
½
½�	½{
½�	½�	½P   P   %
½
½{
½2
½Q
½C
½'
½U
½
½�	½�	½
½h
½
½P
½L
½/
½�
½
½
½P   P   �	½�	½
½�	½)
½�	½'
½
½�	½
½z	½
½
½!
½'
½�	½Y
½�	½�	½�	½P   P   �	½�	½�
½�	½�	½
½�	½3
½
½u
½�	½�	½n
½�	½5
½�	½
½�	½�	½�
½P   P   �	½�	½
½�	½�	½
½�	½�	½~	½�	½%
½
½
½�	½�	½�	½�	½
½
½�	½P   P   �	½
½�	½�	½�	½
½�	½!
½�	½;
½
½0
½2
½�	½1
½�	½
½�	½
½�	½P   P   Y
½

½�	½$
½*
½
½�	½
½�	½[
½:
½�	½f
½�	½8
½[
½�	½
½�	½
½P   P   �	½�	½ 
½
½�	½�	½x	½�	½�	½e
½�	½�	½
½�	½�	½�	½[
½�	½�	½�	½P   P   '
½<
½�	½�	½�	½
½(
½C
½v	½5
½:
½�	½_
½�	½�
½�	½8
½1
½�	½5
½P   P   !
½�	½%
½K
½z
½[
½�	½
½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½P   P   
½�	½�	½9
½3
½�	½�	½�	½
½{
½
½B
½B
½�	½_
½
½f
½2
½
½n
½P   P   
½�	½�	½�	½�	½�	½�	½�	½
½�	½�	½�	½B
½�	½�	½�	½�	½0
½
½�	½P   P   z	½>
½�	½%
½4
½
½�	½
½�	½D
½�	½�	½
½�	½:
½�	½:
½
½%
½�	½P   P   
½F
½�	½�	½ 
½�	½�	½D
½�	½|	½D
½�	½{
½�	½5
½e
½[
½;
½�	½u
½P   P   �	½�	½�	½�	½R
½�	½,
½�	½
½�	½�	½
½
½�	½v	½�	½�	½�	½~	½
½P   P   
½�	½�	½&
½!
½�	½
½�	½�	½D
½
½�	½�	½
½C
½�	½
½!
½�	½3
½P   P   '
½
½�	½�	½
½�	½
½
½,
½�	½�	½�	½�	½�	½(
½x	½�	½�	½�	½�	½P   P   �	½
½@
½0
½�	½�	½�	½�	½�	½�	½
½�	½�	½[
½
½�	½
½
½
½
½P   P   )
½�	½�	½X
½
½�	½
½!
½R
½ 
½4
½�	½3
½z
½�	½�	½*
½�	½�	½�	½P   P   �	½%
½�	½
½X
½0
½�	½&
½�	½�	½%
½�	½9
½K
½�	½
½$
½�	½�	½�	½P   P   
½�	½�	½�	½�	½@
½�	½�	½�	½�	½�	½�	½�	½%
½�	½ 
½�	½�	½
½�
½P   P   �	½�	½�	½%
½�	½
½
½�	½�	½F
½>
½�	½�	½�	½<
½�	½

½
½�	½�	½P   P   �½�	½
½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½{	½�	½!
½�	½
½�	½P   P   �	½
½z	½t	½
½�	½�	½�	½ 
½�	½�	½�	½�	½�	½�	½
½�	½�	½{	½�	½P   P   
½P
½�	½�	½6
½�	½
½
½�	½�	½�	½�
½x	½�	½�	½
½�	½�	½q
½{	½P   P   �	½�	½�	½�	½�	½�	½�	½�	½U	½�	½i	½v	½s	½U	½�	½a	½�	½�	½�	½�	½P   P   !
½l	½�	½t	½�	½�	½

½�	½�	½�	½�	½�	½�	½$
½�	½�	½�	½�	½�	½�	½P   P   �	½{	½?
½%
½�	½�	½�	½
½g	½�	½'	½ 
½�	½�	½�	½@	½�	½a	½
½
½P   P   {	½�	½�	½�	½�	½�	½{	½
½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½P   P   �	½�	½w	½-	½b	½�	½�	½�	½�	½�	½K	½
½�	½�	½�	½�	½$
½U	½�	½�	½P   P   �	½%
½
½�	½
½�	½
½-
½�	½�	½y	½�	½�	½�	½�	½�	½�	½s	½x	½�	½P   P   �	½�	½
½�	½�	½�	½�	½�	½�	½�	½�	½�
½�	½
½�	½ 
½�	½v	½�
½�	½P   P   �	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½y	½K	½�	½'	½�	½i	½�	½�	½P   P   �	½�	½�	½
½�	½�	½�	½�	½	
½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½P   P   �	½�	½�	½	
½�	½�	½F
½�	½�	½	
½�	½�	½�	½�	½�	½g	½�	½U	½�	½ 
½P   P   �	½P
½
½�	½�	½�	½}	½S	½�	½�	½�	½�	½-
½�	½
½
½�	½�	½
½�	½P   P   �	½�	½�	½�	½�	½
½
½}	½F
½�	½�	½�	½
½�	½{	½�	½

½�	½
½�	½P   P   �	½�	½�	½�	½�	½�	½
½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½P   P   �	½�	½�	½N	½�	½�	½�	½�	½�	½�	½�	½�	½
½b	½�	½�	½�	½�	½6
½

½P   P   �	½�	½)
½�	½N	½�	½�	½�	½	
½
½�	½�	½�	½-	½�	½%
½t	½�	½�	½t	½P   P   
½�	½�	½)
½�	½�	½�	½
½�	½�	½�	½
½
½w	½�	½?
½�	½�	½�	½z	½P   P   �	½I
½�	½�	½�	½�	½�	½P
½�	½�	½�	½�	½%
½�	½�	½{	½l	½�	½P
½
½P   P   a
½�	½I	½�	½Y	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½�	½r	½�	½o	½�	½P   P   �	½�	½7	½�	½`	½;	½p	½
	½u	½|	½a	½n	½w	½b	½ 	½�	½B	½H	½�	½	½P   P   o	½	½(	½�	½�	½p	½�	½R	½�	½	
½�	½?	½�	½ 
½�	½L	½�	½m	½�	½�	½P   P   �	½�	½�	½�	½T	½p	½�	½�	½�	½w	½
½�	½�	½
½l	½�	½�	½
½m	½H	½P   P   r	½�	½
½�	½K	½F	½�	½�	½�	½�	½D	½�	½_	½�	½S	½~	½�	½�	½�	½B	½P   P   �	½�	½	½�½�	½�	½m	½H	½�	½|	½�	½�	½�	½~	½�	½�	½~	½�	½L	½�	½P   P   �	½�	½!
½�	½-
½�	½�	½	½�	½k	½Y	½�	½�½�	½	½�	½S	½l	½�	½ 	½P   P   �	½�	½}	½�	½�	½{	½�	½�	½R	½&
½
½�	½�	½
½�	½~	½�	½
½ 
½b	½P   P   �	½|	½b	½�	½�	½�	½|	½z	½�	½|	½�	½�	½X	½�	½�½�	½_	½�	½�	½w	½P   P   �	½�	½K	½�	½�	½�	½�	½.	½�	½�	½l	½8	½�	½�	½�	½�	½�	½�	½?	½n	½P   P   �	½D	½�	½V	½�	½�	½�	½c	½�	½?	½�	½l	½�	½
½Y	½�	½D	½
½�	½a	½P   P   �	½@	½�	½�	½k	½O	½P	½b	½�	½�	½?	½�	½|	½&
½k	½|	½�	½w	½	
½|	½P   P   �	½v	½�	½�	½n	½�	½S	½�	½z	½�	½�	½�	½�	½R	½�	½�	½�	½�	½�	½u	½P   P   �	½�	½G	½^	½a	½�	½�	½�	½�	½b	½c	½.	½z	½�	½	½H	½�	½�	½R	½
	½P   P   �	½�	½Q	½�	½�	½Z	½8	½�	½S	½P	½�	½�	½|	½�	½�	½m	½�	½�	½�	½p	½P   P   �	½�	½�	½�	½�	½�	½Z	½�	½�	½O	½�	½�	½�	½{	½�	½�	½F	½p	½p	½;	½P   P   Y	½�	½
½�	½�	½�	½�	½a	½n	½k	½�	½�	½�	½�	½-
½�	½K	½T	½�	½`	½P   P   �	½�	½	½u	½�	½�	½�	½^	½�	½�	½V	½�	½�	½�	½�	½�½�	½�	½�	½�	½P   P   I	½�	½�	½	½
½�	½Q	½G	½�	½�	½�	½K	½b	½}	½!
½	½
½�	½(	½7	½P   P   �	½	½�	½�	½�	½�	½�	½�	½v	½@	½D	½�	½|	½�	½�	½�	½�	½�	½	½�	½P   P   �½D	½�	½&	½�	½=	½�	½�	½q	½I	½;	½_	½l	½�	½w	½B	½�	½	½�	½H	½P   P   H	½:	½�	½_	½W	½�	½�	½�	½�	½z	½o	½d	½q	½�	½�	½�	½�	½	½W	½�	½P   P   �	½�	½�	½R	½�½�	½0	½�	½I	½�½k	½]	½q	½�½A	½�	½%	½�	½�½W	½P   P   	½	½N	½	½`	½�	½)	½�½�	½*	½N	½�	½�	½H	½(	½�	½�½;	½�	½	½P   P   �	½�	½�	½m	½�	½�	½*	½	½	½J	½>	½�½^	½�½E	½L	½	½�½%	½�	½P   P   B	½u	½D	½H	½q	½)	½�	½�	½�	½N	½�	½.	½�	½�	½1	½�	½L	½�	½�	½�	½P   P   w	½�½ 	½�	½"	½�½�	½�	½H	½4	½9	½/	½R	½*	½J	½1	½E	½(	½A	½�	½P   P   �	½q	½E	½z	½P	½9	½|	½y	½�	½�½I	½�½�	½*	½*	½�	½�½H	½�½�	½P   P   l	½�½�	½b	½	½�	½�	½�½�	½x	½r	½�	½^	½�	½R	½�	½^	½�	½q	½q	½P   P   _	½�	½�	½}	½	½	½`	½�	½�	½6	½d	½b	½�	½�½/	½.	½�½�	½]	½d	½P   P   ;	½b	½�	½�	½X	½6	½c	½�	½�	½h	½^	½d	½r	½I	½9	½�	½>	½N	½k	½o	½P   P   I	½t	½	½�½�	½�	½�	½�	½�½	½h	½6	½x	½�½4	½N	½J	½*	½�½z	½P   P   q	½�	½�	½�½m	½D	½
	½B	½s	½�½�	½�	½�	½�	½H	½�	½	½�	½I	½�	½P   P   �	½�½�	½�	½�	½D	½c	½m	½B	½�	½�	½�	½�½y	½�	½�	½	½�½�	½�	½P   P   �	½g	½�	½y	½Q	½�	½	½c	½
	½�	½c	½`	½�	½|	½�	½�	½*	½)	½0	½�	½P   P   =	½�½=	½f	½	½N	½�	½D	½D	½�	½6	½	½�	½9	½�½)	½�	½�	½�	½�	½P   P   �	½[	½	½k	½"	½	½Q	½�	½m	½�	½X	½	½	½P	½"	½q	½�	½`	½�½W	½P   P   &	½{	½]	½a	½k	½f	½y	½�	½�½�½�	½}	½b	½z	½�	½H	½m	½	½R	½_	½P   P   �	½=	½v	½]	½	½=	½�	½�	½�	½	½�	½�	½�	½E	½ 	½D	½�	½N	½�	½�	½P   P   D	½�	½=	½{	½[	½�½g	½�½�	½t	½b	½�	½�½q	½�½u	½�	½	½�	½:	½P   P   �	½	½		½	½�½�½�½�½	½{½=	½�½�½�½�½	½�½�½!	½	½P   P   	½�½�½	½M	½�½	½�½:	½@	½q	½Q	½8	½S	½�½�½�½�	½�½�½P   P   !	½i	½:	½�½b	½	½	½
	½	½8	½	½�½	½-	½	½	½	½�½1	½�½P   P   �½	½	½�½l	½�½/	½�	½�½�	½>	½�½	½D	½�	½�½�	½5	½�½�	½P   P   �½	½�½�½	½�½	½�	½�½�½�	½	½'	½�½�	½�½�½�	½	½�½P   P   	½t	½S	½	½T	½�½	½	½�½�½�½ 	½	½4	½	½�½�½�½	½�½P   P   �½t	½�½`	½	½�	½�½�½	½�	½�	½	½�	½�½�	½	½�	½�	½	½�½P   P   �½J	½W	½ 	½�½V	½U	½{½^	½
	½J	½	½ 	½�½�½4	½�½D	½-	½S	½P   P   �½]	½'	½	½P	½@	½	½N	½	½<	½%	½�½0	½ 	½�	½	½'	½	½	½8	½P   P   �½	½	½	½�	½|	½�½6	½	½�½V	½�½�½	½	½ 	½	½�½�½Q	½P   P   =	½H	½�½�½�½
	½�½�½�½U	½S	½V	½%	½J	½�	½�½�	½>	½	½q	½P   P   {½d	½B	½d	½�½<	½9	½�½c	½c	½U	½�½<	½
	½�	½�½�½�	½8	½@	½P   P   	½#	½�½^	½I	½�½	½�½U	½c	½�½	½	½^	½	½�½�½�½	½:	½P   P   �½>	½�½�½	½�½2	½I	½�½�½�½6	½N	½{½�½	½�	½�	½
	½�½P   P   �½<	½H	½	½�½)	½�	½2	½	½9	½�½�½	½U	½�½	½	½/	½	½	½P   P   �½�	½E	½�½|	½=	½)	½�½�½<	½
	½|	½@	½V	½�	½�½�½�½	½�½P   P   �½O	½	½�½x	½|	½�½	½I	½�½�½�	½P	½�½	½T	½	½l	½b	½M	½P   P   	½�½t	½@	½�½�½	½�½^	½d	½�½	½	½ 	½`	½	½�½�½�½	½P   P   		½	½�½t	½	½E	½H	½�½�½B	½�½	½'	½W	½�½S	½�½	½:	½�½P   P   	½~	½	½�½O	½�	½<	½>	½#	½d	½H	½	½]	½J	½t	½t	½	½	½i	½�½P   P   [	½�½�½3	½�½	½	½	½'	½�½�½	½	½	½&	½1	½�½!	½�½�½P   P   �½�½,	½	½�½�½7	½�½�½�½�½�½�½�½�½(	½�½�½	½(	½P   P   �½<½�½�½�½�½	½�½�½	½�½�½	½	½�½�½	½�½�½	½P   P   !	½E	½/	½&	½�½�½�½�½�½t½f½�½	½l½y½½�½�½�½�½P   P   �½ 	½�½	½�½�½	½�½U	½(	½�½B	½	½"	½�½,	½Q	½�½	½�½P   P   1	½�½q½�½�½&	½R	½�½u½'	½�½�½T½|½�½�½,	½½�½(	½P   P   &	½�½�½�½�½�½	½�½	½�½�½�½�½#	½�½�½�½y½�½�½P   P   	½�½�½1	½	½�½�½	½�½�½y½,	½`½	½#	½|½"	½l½	½�½P   P   	½2	½W½�½�½�½;½8	½�½�½	½�½7	½`½�½T½	½	½	½�½P   P   	½	½�½	½�½�½�½�½	½#	½�½�½�½,	½�½�½B	½�½�½�½P   P   �½�½�½A	½	½�½/	½L	½m½�½�½�½	½y½�½�½�½f½�½�½P   P   �½�½�½�½�½�½�½�½�½�½�½#	½�½�½�½'	½(	½t½	½�½P   P   '	½/	½�½�½�½2	½�½,	½�½�½m½	½�½�½	½u½U	½�½�½�½P   P   	½	½�½L	½�½3	½�½�½,	½�½L	½�½8	½	½�½�½�½�½�½�½P   P   	½�½w½	½	½�½�½�½�½�½/	½�½;½�½	½R	½	½�½	½7	½P   P   	½�½�½�½�½�½�½3	½2	½�½�½�½�½�½�½&	½�½�½�½�½P   P   �½�½�½+	½�½�½	½�½�½�½	½�½�½	½�½�½�½�½�½�½P   P   3	½	½�½�½+	½�½	½L	½�½�½A	½	½�½1	½�½�½	½&	½�½	½P   P   �½6	½	½�½�½�½w½�½�½�½�½�½W½�½�½q½�½/	½�½,	½P   P   �½@½6	½	½�½�½�½	½/	½�½�½	½2	½�½�½�½ 	½E	½<½�½P   P   �½�½�½9½�½s½g½�½G½�½r½�½G½�½g½s½�½:½�½�½P   P   �½�½�½T½w½�½½~½½^½�½k½k½½u½½�½x½N½�½P   P   �½�½�½:½e½�½�½�½�½�½�½�½�½�½	½�½�½�½c½N½P   P   :½T½:½J½�½�½�½a½�½�½~½n½l½�½�½�½h½�½�½x½P   P   �½w½e½�½�½�½�½d½�½~½w½�½C½�½�½q½�½h½�½�½P   P   s½�½�½�½�½�½3½�½�½a½�½�½�½�½�½�½q½�½�½½P   P   g½½�½�½�½7½;½f½�½�½�½�½5½�½½�½�½�½	½u½P   P   �½�½�½a½d½�½h½	½?½�½�½�½�½�½�½�½�½�½�½½P   P   G½½�½�½�½�½�½=½½Q½�½a½l½�½5½�½C½l½�½k½P   P   �½\½�½�½�½d½�½�½N½>	½y½�½a½�½�½�½�½n½�½k½P   P   r½�½�½z½u½�½�½�½�½w½$½y½�½�½�½�½w½~½�½�½P   P   �½j½�½n½�½�½�½�½`½�½w½>	½Q½�½�½a½~½�½�½^½P   P   G½h½�½l½D½�½5½�½n½`½�½N½½?½�½�½�½�½�½½P   P   �½½�½}½�½�½�½�½�½�½�½�½=½	½f½�½d½a½�½~½P   P   g½x½	½�½}½�½½�½5½�½�½�½�½h½;½3½�½�½�½½P   P   s½½�½�½s½�½�½�½�½�½�½d½�½�½7½�½�½�½�½�½P   P   �½�½�½g½�½s½}½�½D½�½u½�½�½d½�½�½�½�½e½w½P   P   9½x½�½�½g½�½�½}½l½n½z½�½�½a½�½�½�½J½:½T½P   P   �½N½c½�½�½�½	½�½�½�½�½�½�½�½�½�½e½:½�½�½P   P   �½�½N½x½�½½x½½h½j½�½\½½�½½�½w½T½�½�½P   P   �½H½ ½�½½�½�½o½�½o½T½K½�½�½�½�½>½�½$½D½P   P   D½9½�½�½�½/½H½½�½�½9½A½�½�½½h½½n½�½�½P   P   $½�½8½�½e½�½½Z½�½>½�½E½�½)½�½J½½�½½�½P   P   �½s½X½�½�½½K½�½
½v½�½`½[½�½�½½�½8½�½n½P   P   >½'½j½L½4½½½�½½2½x½#½½&½q½½4½�½½½P   P   �½9½$½½"½�½l½W½?½½/½$½�½�½½S½½½J½h½P   P   �½�½}½½�½�½y½½�½]½�½%½-½½:½½q½�½�½½P   P   �½f½½�½½ ½I½�½�½^½�½½�½½½�½&½�½)½�½P   P   �½½d½�½�½�½~½N½f½{½�½Z½>½�½-½�½½[½�½�½P   P   K½/½�½�½�½�½�½M½%½�½@½a½Z½½%½$½#½`½E½A½P   P   T½L½\½�½2½+½(½�½�½2½,½@½�½�½�½/½x½�½�½9½P   P   o½$½)½k½�½A½N½�½^½½2½�½{½^½]½½2½v½>½�½P   P   �½.½q½r½�½�½`½�½�½^½�½%½f½�½�½?½½
½�½�½P   P   o½8½u½�½�½�½�½x½�½�½�½M½N½�½½W½�½�½Z½½P   P   �½f½`½�½;½U½0½�½`½N½(½�½~½I½y½l½½K½½H½P   P   �½�½½�½�½½U½�½�½A½+½�½�½ ½�½�½½½�½/½P   P   ½5½�½½�½�½;½�½�½�½2½�½�½½�½"½4½�½e½�½P   P   �½T½½½½�½�½�½r½k½�½�½�½�½½½L½�½�½�½P   P    ½s½C½½�½½`½u½q½)½\½�½d½½}½$½j½X½8½�½P   P   H½�½s½T½5½�½f½8½.½$½L½/½½f½�½9½'½s½�½9½P   P   c½�½�½�½�½�½�½b½�½�½½T½�½}½�½�½�½�½�½�½P   P   �½�½D½�½�½L½J½#½4½�½#½?½�½½½g½(½�½�½Y½P   P   �½�½½�½�½.½�½/½½�½�½½�½�½$½½�½O½�½�½P   P   �½�½�½�½�½Z½9½�½�½�½�½=½8½�½�½�½�½½O½�½P   P   �½(½;½F½�½-½�½�½(½t½�½�½#½�½�½U½P½�½�½(½P   P   �½�½�½�½�½�½Y½.½½V½�½½�½�½½½U½�½½g½P   P   �½�½�½½�½�½�½-½�½�½�½½Y½½t½½�½�½$½½P   P   }½�½�½|½�½�½�½T½%½½�½�½�½"½½�½�½�½�½½P   P   �½½�½�½�½�½�½8½�½�½�½<½/½�½Y½�½#½8½�½�½P   P   T½½½j½�½�½�½�½½a½0½>½<½�½½½�½=½½?½P   P   ½J½�½½�½z½k½#½�½0½-½0½�½�½�½�½�½�½�½#½P   P   �½+½�½�½�½�½�½�½�½�½0½a½�½½�½V½t½�½�½�½P   P   �½½�½�½�½�½�½�½½�½�½½�½%½�½½(½�½½4½P   P   b½-½½½�½½�½�½�½�½#½�½8½T½-½.½�½�½/½#½P   P   �½�½�½o½�½�½�½�½�½�½k½�½�½�½�½Y½�½9½�½J½P   P   �½�½�½�½�½b½�½½�½�½z½�½�½�½�½�½-½Z½.½L½P   P   �½�½�½~½�½�½�½�½�½�½�½�½�½�½�½�½�½�½�½�½P   P   �½k½�½½~½�½o½½�½�½½j½�½|½½�½F½�½�½�½P   P   �½�½
½�½�½�½�½½�½�½�½½�½�½�½�½;½�½½D½P   P   �½q½�½k½�½�½�½-½½+½J½½½�½�½�½(½�½�½�½P   P   ½�½½]½�½�½�½�½�½�½�½�½�½�½�½�½�½n½�½�½P   P   �½�½�½c½�½�½½�½C½�½�½�½�½A½�½"½�½�½�½�½P   P   �½/½�½�½�½�½H½�½�½�½½E½½�½�½�½a½�½�½�½P   P   n½�½�½\½�½�½�½�½�½�½�½B½9½�½�½�½�½�½�½�½P   P   �½�½½�½ ½�½j½�½[½a½�½½�½½�½W½h½�½a½�½P   P   �½½�½�½½q½½�½�½\½|½�½�½�½�½�½W½�½�½"½P   P   �½�½s½k½m½�½�½�½�½�½�½�½O½�½Y½�½�½�½�½�½P   P   �½½�½?½J½�½½�½4½�½�½ ½�½�½�½�½½�½�½A½P   P   �½�½�½
½X½½�½�½�½�½ ½<½�½�½O½�½�½9½½�½P   P   �½�½�½n½�½�½x½�½�½½�½L½<½ ½�½�½½B½E½�½P   P   �½�½�½�½�½(½~½�½�½�½�½�½ ½�½�½|½�½�½½�½P   P   �½�½�½�½½v½w½½�½�½�½½�½�½�½\½a½�½�½�½P   P   �½�½�½�½�½�½�½�½�½�½�½�½�½4½�½�½[½�½�½C½P   P   �½�½½�½½�½q½q½�½½�½�½�½�½�½�½�½�½�½�½P   P   �½½�½l½�½y½�½q½�½w½~½x½�½½�½½j½�½H½½P   P   �½�½�½½�½ ½y½�½�½v½(½�½½�½�½q½�½�½�½�½P   P   �½½h½?½S½�½�½½�½½�½�½X½J½m½½ ½�½�½�½P   P   ]½�½�½~½?½½l½�½�½�½�½n½
½?½k½�½�½\½�½c½P   P   ½�½�½�½h½�½�½½�½�½�½�½�½�½s½�½½�½�½�½P   P   �½½�½�½½�½½�½�½�½�½�½�½½�½½�½�½/½�½P   P   ½K½ ½b½%½G½[½`½Q½�½d½�½J½=½s½_½½b½�½I½P   P   I½g½�½>½T½A½�½`½2½?½�½�½*½S½e½y½O½X½e½�½P   P   �½�½�½u½�½�½�½/½½ ½F½�½U½�½½9½�½�½�½e½P   P   b½�½�½z½@½�½6½t½I½D½	½r½h½½=½O½�½'½�½X½P   P   ½½`½½�½j½�½½X½g½W½½!½½W½|½5½�½�½O½P   P   _½�½&½%½�½a½m½-½5½v½�½½�½�½½k½|½O½9½y½P   P   s½#½S½�½T½ ½i½g½0½C½S½½½~½�½½W½=½½e½P   P   =½�½½R½R½�½�½R½0½�½½½�½m½~½�½½½�½S½P   P   J½'½E½g½�½t½H½½^½@½^½f½,½�½½�½!½h½U½*½P   P   �½.½�½,½=½/½½�½.½�½�½|½f½½½½½r½�½�½P   P   d½½G½�½�½�½½�½C½ ½m½�½^½½S½�½W½	½F½�½P   P   �½"½�½4½�½�½x½�½;½�½ ½�½@½�½C½v½g½D½ ½?½P   P   Q½)½F½1½½H½�½:½	½;½C½.½^½0½0½5½X½I½½2½P   P   `½½�½�½�½/½�½�½:½�½�½�½½R½g½-½½t½/½`½P   P   [½�½F½!½½q½�½�½�½x½½½H½�½i½m½�½6½�½�½P   P   G½G½½w½1½�½q½/½H½�½�½/½t½�½ ½a½j½�½�½A½P   P   %½�½9½P½�½1½½�½½�½�½=½�½R½T½�½�½@½�½T½P   P   b½�½#½�½P½w½!½�½1½4½�½,½g½R½�½%½½z½u½>½P   P    ½�½w½#½9½½F½�½F½�½G½�½E½½S½&½`½�½�½�½P   P   K½�½�½�½�½G½�½½)½"½½.½'½�½#½�½½�½�½g½P   P   ½½,½½C½�½�½�½�½�½�½�½�½�½�½�½ ½�½;½½P   P   ½/½r½�½�½�½�½�½C½�½½�½�½o½�½�½�½�½�½k½P   P   ;½�½½�½�½`½½�½:½8½�½½�½:½½�½½J½�½�½P   P   �½�½�½½�½F½�½M½½�½�½*½&½�½�½½n½�½J½�½P   P    ½*½S½½�½�½�½�½(½�½½�½�½�½�½�½�½n½½�½P   P   �½�½�½�½½½�½�½�½�½�½ ½�½�½"½�½�½½�½�½P   P   �½½ ½�½'½½�½�½:½½�½½g½�½7½"½�½�½½�½P   P   �½½;½�½�½.½*½�½K½½�½�½�½r½�½�½�½�½:½o½P   P   �½!½½s½�½�½½�½�½�½�½&½�½�½g½�½�½&½�½�½P   P   �½�½�½½½½�½½�½�½�½½&½�½½ ½�½*½½�½P   P   �½�½�½�½�½F½�½i½�½½�½�½�½�½�½�½½�½�½½P   P   �½½�½�½½ ½½7½�½�½½�½�½½½�½�½�½8½�½P   P   �½�½�½�½�½�½�½�½�½�½�½�½�½K½:½�½(½½:½C½P   P   �½�½½s½C½�½�½½�½7½i½½�½�½�½�½�½M½�½�½P   P   �½½½�½�½�½½�½�½½�½�½½*½�½�½�½�½½�½P   P   �½:½5½½½`½�½�½�½ ½F½½�½.½½½�½F½`½�½P   P   C½½½�½�½½�½C½�½½�½½�½�½'½½�½�½�½�½P   P   ½�½�½�½�½½�½s½�½�½�½½s½�½�½�½½½�½�½P   P   ,½�½�½�½½5½½½�½�½�½�½½;½ ½�½S½�½½r½P   P   ½�½�½�½½:½½�½�½½�½�½!½½½�½*½�½�½/½P   P   (½d½k½}½�½o½�½�½�½�½	½�½�½�½�½�½�½l½�½e½P   P   e½m½½�½�½3½�½|½½�½�½�½{½.½�½�½V½�½y½½P   P   �½½�½z½X½�½R½�½I½u½z½½m½�½½�½H½�½y½y½P   P   l½Y½c½o½�½�½½�½�½½�½'½2½�½.½�½�½�½�½�½P   P   �½@½W½5½�½X½&½½�½+½�½�½�½�½�½R½�½�½H½V½P   P   �½�½�½�½�½�½�½�½{½b½�½-½]½L½P½�½R½�½�½�½P   P   �½½9½.½8½½�½�½-½T½�½?½�½�½�½P½�½.½½�½P   P   �½�½{½�½�½�½�½�½½y½�½�½d½t½�½L½�½�½�½.½P   P   �½�½½j½l½g½½}½�½�½k½=½�½d½�½]½�½2½m½{½P   P   �½½½�½�½�½�½8½	½z½�½½=½�½?½-½�½'½½�½P   P   	½'½�½�½�½l½�½x½�½;½ ½�½k½�½�½�½�½�½z½�½P   P   �½D½�½�½?½w½i½_½�½�½;½z½�½y½T½b½+½½u½�½P   P   �½�½�½�½�½�½�½�½�½�½�½	½�½½-½{½�½�½I½½P   P   �½�½1½�½]½g½8½M½�½_½x½8½}½�½�½�½½�½�½|½P   P   �½�½½�½�½e½½8½�½i½�½�½½�½�½�½&½½R½�½P   P   o½½|½i½�½y½e½g½�½w½l½�½g½�½½�½X½�½�½3½P   P   �½�½<½�½v½�½�½]½�½?½�½�½l½�½8½�½�½�½X½�½P   P   }½½�½3½�½i½�½�½�½�½�½�½j½�½.½�½5½o½z½�½P   P   k½R½�½�½<½|½½1½�½�½�½½½{½9½�½W½c½�½½P   P   d½N½R½½�½½�½�½�½D½'½½�½�½½�½@½Y½½m½P   P   }½½�½,½�½½½�½½½�½�½½�½
½½�½%½�½½P   P   ½½½�½)½F½G½½d½�½�½�½½Q½ ½:½K½+½v½½P   P   �½�½�½u½�½�½½�½C½(½�½�½g½B½5½�½½�½�½v½P   P   %½�½�½½B½�½ ½�½½A½�½#½4½�½E½½�½B½�½+½P   P   �½�½½�½�½=½½ ½f½b½(½�½}½�½½q½}½�½½K½P   P   ½8½_½Z½J½½=½�½�½�½{½½)½�½½v½q½½�½:½P   P   
½½=½4½0½½½½:½]½�½�½5½,½_½½½E½5½ ½P   P   �½�½ ½@½K½;½�½�½P½;½�½!½!½.½,½�½�½�½B½Q½P   P   ½�½c½p½�½P½W½�½%½½o½I½!½!½5½)½}½4½g½½P   P   �½
½$½�½T½u½½0½½�½�½s½I½!½�½½�½#½�½�½P   P   �½S½:½�½½l½�½w½-½X½�½�½o½�½�½{½(½�½�½�½P   P   ½T½C½�½�½�½½�½�½C½X½�½½;½]½�½b½A½(½�½P   P   ½�½<½�½#½½!½½�½�½-½½%½P½:½�½f½½C½d½P   P   �½�½9½u½�½½'½½½�½w½0½�½�½½�½ ½�½�½½P   P   ½½V½�½½
½!½'½!½½�½½W½�½½=½½ ½½G½P   P   ½�½(½i½i½T½
½½½�½l½u½P½;½½½=½�½�½F½P   P   �½I½F½@½�½i½½�½#½�½½T½�½K½0½J½�½B½�½)½P   P   ,½�½O½5½@½i½�½u½�½�½�½�½p½@½4½Z½�½½u½�½P   P   �½�½½O½F½(½V½9½<½C½:½$½c½ ½=½_½½�½�½½P   P   ½�½�½�½I½�½½�½�½T½S½
½�½�½½8½�½�½�½½P   P   +½�½�½�½�½�½�½�½�½�½�½�½�½�½�½y½�½�½�½�½P   P   �½�½Z½Q½�½�½d½�½�½�½S½f½�½�½�½�½�½r½R½\½P   P   �½�½�½U½�½�½�½�½�½I½�½�½�½m½�½�½�½�½�½R½P   P   �½�½�½�½�½�½�½�½�½�½�½r½v½�½�½�½�½�½�½r½P   P   �½�½;½�½�½�½�½�½�½�½g½�½g½�½�½{½�½�½�½�½P   P   y½�½[½J½�½�½r½x½�½�½½!½�½�½�½½{½�½�½�½P   P   �½E½�½�½�½%½�½�½�½�½t½�½�½\½�½�½�½�½�½�½P   P   �½�½6½½1½R½�½�½�½a½�½�½�½�½\½�½�½�½m½�½P   P   �½�½�½�½½�½�½�½�½�½�½�½1½�½�½�½g½v½�½�½P   P   �½0½�½P½�½½k½�½8½�½o½�½�½�½�½!½�½r½�½f½P   P   �½�½�½n½�½/½�½s½�½�½�½o½�½�½t½½g½�½�½S½P   P   �½�½O½�½�½�½�½½�½M½�½�½�½a½�½�½�½�½I½�½P   P   �½½�½�½�½�½]½�½�½�½�½8½�½�½�½�½�½�½�½�½P   P   �½½�½a½�½�½�½�½�½½s½�½�½�½�½x½�½�½�½�½P   P   �½�½�½Q½�½�½>½�½]½�½�½k½�½�½�½r½�½�½�½d½P   P   �½ ½D½�½½�½�½�½�½�½/½½�½R½%½�½�½�½�½�½P   P   �½�½�½&½�½½�½�½�½�½�½�½½1½�½�½�½�½�½�½P   P   �½½M½�½&½�½Q½a½�½�½n½P½�½½�½J½�½�½U½Q½P   P   �½�½&½M½�½D½�½�½�½O½�½�½�½6½�½[½;½�½�½Z½P   P   �½�½�½½�½ ½�½½½�½�½0½�½�½E½�½�½�½�½�½P   