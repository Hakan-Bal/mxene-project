H   e�ݯ>@K����c�a�ӄ�3?����B��9�7 @�D�߅�3��w��rc?֐��oV�=xU=-�E@H            �         P   ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ%�Ͻ8�Ͻ��Ͻ��Ͻ��ϽU�Ͻ��Ͻ��Ͻl�Ͻ��Ͻ3�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ=�Ͻ��Ͻ1�Ͻo�Ͻ��Ͻ��Ͻ��Ͻ9�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ~�ϽP�Ͻ"�Ͻ(�Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻ�Ͻh�Ͻ��Ͻ��Ͻ��Ͻ@�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ1�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ(�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ3�Ͻ��Ͻ��Ͻ��Ͻ�Ͻl�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻc�Ͻ��Ͻ"�ϽP   P   ��ϽM�ϽY�Ͻ*�Ͻ��Ͻ/�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ8�Ͻ��Ͻ��ϽB�Ͻ��Ͻ��Ͻ��ϽP�ϽP   P   3�Ͻ��Ͻ��Ͻ��Ͻc�Ͻ8�Ͻj�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ}�ϽB�Ͻ�Ͻ��Ͻ~�ϽP   P   ��Ͻ��Ͻr�Ͻ �Ͻ��Ͻ��Ͻ.�Ͻ��Ͻ\�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   l�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻt�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ1�Ͻ��ϽP   P   ��Ͻ?�Ͻ��Ͻ��ϽM�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ<�Ͻ{�ϽU�Ͻ��Ͻ��Ͻ��Ͻ8�Ͻ��Ͻ��Ͻ��ϽP   P   ��ϽS�Ͻ$�Ͻ��Ͻ��Ͻ	�Ͻ��Ͻ`�Ͻ=�Ͻ��Ͻ��Ͻ��Ͻ{�Ͻ��Ͻ��Ͻ��Ͻ��Ͻl�Ͻ��Ͻ��ϽP   P   U�Ͻa�Ͻ��Ͻ8�Ͻ�Ͻ��Ͻ#�Ͻ�Ͻ��Ͻc�Ͻ��Ͻ��Ͻ<�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ9�ϽP   P   ��Ͻv�Ͻ��Ͻ��ϽP�Ͻ��Ͻ��Ͻt�Ͻ��Ͻ��Ͻc�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ~�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ=�Ͻ��Ͻ��Ͻ\�Ͻ��Ͻ��Ͻ��Ͻ@�Ͻ��ϽP   P   ��Ͻ��Ͻ�Ͻ+�Ͻr�Ͻu�Ͻ��Ͻ��Ͻ��Ͻt�Ͻ�Ͻ`�Ͻ��Ͻt�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   8�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ#�Ͻ��Ͻ��Ͻ��Ͻ.�Ͻj�Ͻ��Ͻ3�Ͻ��Ͻo�ϽP   P   %�Ͻ��Ͻ��ϽY�Ͻ��Ͻ��Ͻ��Ͻu�Ͻ��Ͻ��Ͻ��Ͻ	�Ͻ��Ͻ��Ͻ��Ͻ8�Ͻ/�Ͻ��Ͻ��Ͻ1�ϽP   P   �Ͻj�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻr�Ͻ�ϽP�Ͻ�Ͻ��ϽM�Ͻ��Ͻ��Ͻc�Ͻ��Ͻ��Ͻh�Ͻ��ϽP   P   ��Ͻ�Ͻ��Ͻ��Ͻ��ϽY�Ͻ��Ͻ+�Ͻ��Ͻ��Ͻ8�Ͻ��Ͻ��Ͻ�Ͻ �Ͻ��Ͻ*�Ͻ��Ͻ�Ͻ=�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ$�Ͻ��Ͻ��Ͻr�Ͻ��ϽY�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ�Ͻ��Ͻ�Ͻj�Ͻ��Ͻ��Ͻ��Ͻ~�Ͻv�Ͻa�ϽS�Ͻ?�Ͻ��Ͻ��Ͻ��ϽM�Ͻ��Ͻ��Ͻ��ϽP   P   }�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽU�Ͻ��Ͻ��Ͻ �Ͻ6�Ͻ��ϽJ�Ͻ��Ͻ|�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽZ�Ͻ��Ͻ��Ͻ��Ͻ%�Ͻ��Ͻ��Ͻ�Ͻ��ϽZ�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ'�Ͻ��Ͻ��Ͻ��Ͻ��Ͻr�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻu�Ͻ��ϽP   P   ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ>�Ͻ�Ͻ��Ͻ��Ͻ��Ͻe�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻl�Ͻ��Ͻ��ϽP   P   ��Ͻ��ϽI�Ͻ��Ͻ��Ͻx�Ͻ&�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   |�ϽC�Ͻ��Ͻ�Ͻ�Ͻ��ϽZ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻv�Ͻ��Ͻ��Ͻ��ϽZ�ϽP   P   ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽB�Ͻ%�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   J�Ͻ �ϽC�Ͻ��Ͻ��Ͻ`�Ͻ��ϽZ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ%�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻq�Ͻ��Ͻv�Ͻ�Ͻ��Ͻ�Ͻh�Ͻ��Ͻ�ϽB�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   6�Ͻ��Ͻn�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ*�Ͻ��Ͻ^�Ͻh�Ͻ��Ͻ��Ͻ��Ͻ��Ͻe�Ͻr�Ͻ��ϽP   P    �Ͻj�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽV�Ͻ0�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ%�ϽP   P   ��Ͻv�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�ϽV�Ͻ*�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ2�Ͻ��Ͻ3�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   U�Ͻ]�Ͻ_�Ͻ��Ͻ��Ͻ0�Ͻ��Ͻ��Ͻ3�Ͻ��Ͻ��Ͻ��Ͻv�ϽZ�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ�Ͻy�Ͻ�Ͻd�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽZ�Ͻ&�Ͻ>�Ͻ'�ϽZ�ϽP   P   ��Ͻ��ϽT�ϽC�Ͻ��Ͻ��Ͻ�Ͻ0�Ͻ2�Ͻ��Ͻ��Ͻ��Ͻq�Ͻ`�Ͻ��Ͻ��Ͻx�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ9�Ͻ�Ͻ��Ͻ�Ͻ��Ͻy�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��ϽC�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻj�Ͻ��Ͻ�ϽT�Ͻ��Ͻ_�Ͻ��Ͻ�Ͻ��Ͻn�Ͻ��ϽC�Ͻ�Ͻ��ϽI�Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ$�Ͻ��Ͻ��Ͻ9�Ͻ��Ͻ��Ͻ]�Ͻ�Ͻv�Ͻj�Ͻ��Ͻ��Ͻ �Ͻ�ϽC�Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   y�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ$�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ�Ͻ��Ͻ-�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻz�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ@�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ6�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ"�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   �Ͻx�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ#�Ͻ�Ͻ�Ͻ2�Ͻ�Ͻ&�Ͻ<�Ͻ�ϽP�Ͻ��Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ!�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ6�Ͻ��Ͻ��Ͻl�Ͻ��Ͻ��Ͻ<�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ.�Ͻ��Ͻ��Ͻl�Ͻ��Ͻ&�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻq�Ͻ�Ͻl�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ
�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ��ϽE�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��ϽB�Ͻ
�Ͻ.�Ͻ��Ͻ��Ͻ2�Ͻ"�Ͻ@�Ͻ��ϽP   P   ��Ͻu�Ͻ��Ͻ
�Ͻ�Ͻx�Ͻ��Ͻ2�Ͻ��Ͻ��Ͻf�Ͻ��Ͻ�Ͻ��Ͻ6�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ|�Ͻ��Ͻv�Ͻ��Ͻ��Ͻb�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��ϽX�Ͻ��Ͻ��ϽK�Ͻ��Ͻ$�Ͻb�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ#�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ!�Ͻ�Ͻ:�Ͻ��Ͻ��Ͻ��Ͻs�Ͻ��Ͻ��Ͻ2�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽK�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ!�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   $�Ͻ��Ͻ.�Ͻy�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻv�Ͻx�Ͻ��Ͻl�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ6�Ͻ��Ͻ-�ϽP   P   �Ͻ�Ͻ��Ͻ��Ͻ��Ͻy�Ͻ��Ͻ:�ϽX�Ͻ|�Ͻ
�Ͻ��Ͻq�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ.�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��ϽE�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   ��Ͻr�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ!�Ͻ��Ͻ��Ͻu�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻx�Ͻ��Ͻz�Ͻ��ϽP   P   ��Ͻ7�Ͻ��Ͻ{�ϽX�Ͻ��Ͻ��ϽW�Ͻ��Ͻ�Ͻ0�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ.�ϽP   P   .�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻy�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ �Ͻ��Ͻ��Ͻ{�Ͻ��Ͻ��Ͻ��Ͻi�Ͻ��Ͻ��Ͻ��Ͻ:�Ͻ��ϽP   P   ��Ͻl�Ͻ��Ͻa�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ}�Ͻ��ϽP�Ͻ��Ͻ��Ͻ��Ͻ��Ͻa�Ͻ��Ͻ��Ͻ��Ͻy�ϽP   P   ��Ͻ��Ͻf�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻv�Ͻm�Ͻ��Ͻi�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�ϽP   P   ��ϽM�Ͻ��Ͻ]�Ͻ��Ͻ��Ͻ'�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻa�Ͻ��Ͻ�ϽP   P   ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽO�Ͻ�Ͻ��Ͻ��Ͻ��Ͻi�Ͻ��ϽP   P   ��Ͻ��Ͻ@�Ͻ�Ͻ=�Ͻ�Ͻ��Ͻ^�Ͻ��Ͻ�Ͻk�Ͻ��Ͻ��Ͻ��ϽO�Ͻ��Ͻi�Ͻ��Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽV�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ.�Ͻ'�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻm�Ͻ��Ͻ��Ͻ��ϽP   P   0�Ͻ�Ͻ��Ͻ<�Ͻ��Ͻx�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽV�Ͻk�Ͻ��Ͻ��Ͻv�ϽP�Ͻ{�Ͻ��ϽP   P   �Ͻ�Ͻ��Ͻb�Ͻ�Ͻ��Ͻ��Ͻ��ϽX�Ͻ��Ͻ�Ͻ'�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��ϽS�ϽJ�Ͻ��Ͻ�Ͻ�Ͻc�ϽX�Ͻ��Ͻ.�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ}�Ͻ��Ͻ��ϽP   P   W�Ͻ��Ͻ��Ͻw�Ͻ��Ͻ(�ϽO�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ^�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ �Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽO�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ'�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ=�Ͻ��Ͻ��Ͻd�Ͻ��Ͻ(�Ͻ��Ͻ��Ͻx�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   X�Ͻp�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��ϽJ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ=�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   {�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻw�ϽS�Ͻb�Ͻ<�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ]�Ͻ��Ͻa�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ=�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ@�Ͻ�Ͻ��Ͻf�Ͻ��Ͻ��Ͻ�ϽP   P   7�Ͻ��Ͻ��Ͻ�Ͻp�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��ϽM�Ͻ��Ͻl�Ͻ��Ͻ��ϽP   P   s�ϽK�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ6�Ͻ��Ͻ��Ͻ��Ͻ<�Ͻ��Ͻ_�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽS�ϽP   P   S�ϽC�ϽH�Ͻ��Ͻ��Ͻ�ϽB�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ|�Ͻ��ϽP�Ͻ��Ͻ��Ͻ��Ͻ?�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻq�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ}�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻq�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ3�Ͻ�Ͻ��Ͻ�ϽU�Ͻ��Ͻ��Ͻd�Ͻ��Ͻ��Ͻ��Ͻ	�Ͻ��Ͻ��ϽP   P   �Ͻ��ϽB�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ)�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽQ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻh�Ͻ��Ͻ��Ͻ��Ͻq�Ͻ3�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   _�Ͻ��Ͻ��Ͻ%�Ͻ7�Ͻ��Ͻ��Ͻ=�Ͻ��Ͻ��Ͻc�Ͻ�Ͻ��Ͻa�Ͻ3�Ͻ��Ͻ�Ͻd�Ͻ}�Ͻ|�ϽP   P   ��ϽM�Ͻ��Ͻ��ϽI�Ͻ��Ͻ|�Ͻr�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻq�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   <�ϽG�Ͻ��Ͻ��Ͻ,�Ͻ�Ͻ��Ͻ\�Ͻn�Ͻi�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ7�Ͻ��Ͻ��Ͻ�Ͻm�Ͻ��Ͻ��Ͻ��Ͻc�Ͻ��Ͻ��Ͻ��ϽU�Ͻ��Ͻ��ϽP   P   ��ϽS�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻm�Ͻi�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ]�Ͻ
�Ͻ�Ͻ��Ͻd�Ͻ��Ͻn�Ͻ��Ͻ��Ͻ�Ͻn�Ͻ��Ͻ��Ͻh�Ͻ�Ͻ��Ͻ��Ͻq�Ͻ��ϽP   P   6�Ͻ}�Ͻ��Ͻ}�Ͻ��Ͻp�Ͻ�Ͻ��Ͻn�Ͻ��Ͻ��Ͻ\�Ͻr�Ͻ=�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ��ϽU�Ͻ��Ͻ��Ͻ��Ͻn�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ|�Ͻ��Ͻ��ϽQ�Ͻ��Ͻ3�Ͻ��ϽB�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ/�Ͻ�Ͻ��Ͻp�Ͻd�Ͻ��Ͻ7�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻ6�Ͻ2�Ͻ/�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ,�ϽI�Ͻ7�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ0�Ͻ��Ͻ��Ͻ6�Ͻ��Ͻ��Ͻ}�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ%�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽU�Ͻ��Ͻ
�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽB�Ͻ��Ͻ��ϽH�ϽP   P   K�Ͻ��Ͻ��Ͻ0�Ͻ��Ͻ��Ͻ��Ͻ}�Ͻ]�ϽS�Ͻ��ϽG�ϽM�Ͻ��Ͻ��Ͻ��Ͻ��Ͻq�Ͻ��ϽC�ϽP   P   ��Ͻ��Ͻ��Ͻ3�Ͻ�Ͻ��Ͻ��Ͻw�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻj�Ͻ��Ͻ��Ͻ�ϽA�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ
�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��ϽX�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻd�Ͻ��ϽP   P   A�Ͻ��Ͻ��Ͻb�Ͻr�Ͻ��Ͻ�Ͻ^�Ͻ��Ͻ��Ͻ��Ͻk�Ͻ��Ͻn�Ͻ��Ͻ��Ͻa�Ͻ��Ͻ��Ͻ��ϽP   P   �ϽX�Ͻ��ϽF�ϽG�Ͻ��Ͻ��Ͻ*�Ͻ��Ͻ��Ͻ��Ͻ��Ͻt�Ͻ��Ͻc�Ͻ��Ͻ��Ͻa�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ\�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻs�Ͻ��Ͻz�Ͻ��Ͻ��Ͻ��Ͻ��Ͻj�Ͻ��Ͻ��Ͻ��Ͻ"�Ͻ��Ͻ��Ͻc�Ͻ��Ͻ��Ͻ��ϽP   P   j�Ͻ��Ͻ��Ͻ.�Ͻ�Ͻ��Ͻ��Ͻv�Ͻ��Ͻ��Ͻx�Ͻw�Ͻ��Ͻ
�Ͻ"�Ͻ��Ͻ��Ͻn�Ͻ��Ͻ��ϽP   P   ��Ͻ �Ͻ��Ͻ{�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻx�Ͻ��Ͻ��Ͻ��Ͻ��Ͻt�Ͻ��Ͻ��Ͻ
�ϽP   P   ��Ͻ��Ͻ%�Ͻd�Ͻe�ϽZ�Ͻb�Ͻ:�Ͻ��Ͻ��Ͻ��Ͻ��Ͻx�Ͻw�Ͻ��Ͻ��Ͻ��Ͻk�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻx�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ[�Ͻj�Ͻ��Ͻ��Ͻe�Ͻa�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻj�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻa�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   w�Ͻ��Ͻ4�Ͻ��Ͻt�Ͻ��ϽP�ϽE�Ͻ��Ͻe�Ͻ��Ͻ:�Ͻ��Ͻv�Ͻ��Ͻ�Ͻ*�Ͻ^�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP�Ͻ��Ͻ��Ͻ��Ͻb�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻp�Ͻd�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽZ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�ϽP   P   �Ͻy�Ͻy�Ͻ(�Ͻ��Ͻd�Ͻ��Ͻt�Ͻ��Ͻj�Ͻ��Ͻe�Ͻ��Ͻ�Ͻz�Ͻ\�ϽG�Ͻr�Ͻ��Ͻ��ϽP   P   3�Ͻy�Ͻ��Ͻ��Ͻ(�Ͻp�Ͻ��Ͻ��Ͻ��Ͻ[�Ͻ��Ͻd�Ͻ{�Ͻ.�Ͻ��Ͻ��ϽF�Ͻb�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻy�Ͻ��Ͻ��Ͻ4�Ͻ��Ͻ��Ͻ��Ͻ%�Ͻ��Ͻ��Ͻs�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻw�Ͻ��Ͻy�Ͻy�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ �Ͻ��Ͻ��Ͻ��ϽX�Ͻ��ϽX�Ͻ��ϽP   P   ��Ͻd�Ͻ��Ͻ��Ͻ��Ͻo�Ͻ��ϽT�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ]�Ͻ#�Ͻ��Ͻ��Ͻ��Ͻ��ϽO�Ͻi�ϽP   P   i�Ͻ��Ͻ��ϽX�Ͻ��Ͻ�Ͻ_�Ͻn�Ͻ��Ͻ��Ͻ��Ͻ_�Ͻ��Ͻ��Ͻ��ϽE�Ͻ#�Ͻ
�Ͻb�Ͻ�ϽP   P   O�ϽT�Ͻq�Ͻd�Ͻ��Ͻ��Ͻ��Ͻq�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ	�Ͻ|�Ͻp�Ͻ��Ͻ��Ͻ��Ͻb�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ7�Ͻ�Ͻz�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ=�Ͻ!�Ͻ��Ͻ
�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ+�Ͻ��Ͻ"�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻz�Ͻ=�Ͻ��Ͻ#�ϽP   P   ��Ͻ��Ͻ^�Ͻ��Ͻ��Ͻ��Ͻ;�Ͻn�Ͻk�Ͻ��Ͻ��Ͻ��Ͻ��Ͻm�Ͻ��Ͻ��Ͻ��Ͻ��Ͻp�ϽE�ϽP   P   ��Ͻ��Ͻ[�Ͻ�Ͻa�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ{�Ͻ��Ͻ��Ͻ��Ͻ|�Ͻ��ϽP   P   #�Ͻ��Ͻ��Ͻs�ϽD�Ͻ��Ͻ��ϽZ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻp�Ͻ��Ͻm�Ͻ��Ͻ��Ͻ	�Ͻ��ϽP   P   ]�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻv�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻc�Ͻ��Ͻ��Ͻw�Ͻ_�ϽN�Ͻ+�ϽO�Ͻ��Ͻ[�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ_�ϽP   P   ��Ͻ��ϽO�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ]�Ͻ��Ͻ��Ͻ[�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��ϽJ�Ͻ��Ͻ_�Ͻ_�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻq�Ͻd�Ͻ��Ͻ��Ͻ��Ͻ'�Ͻ��Ͻ��Ͻ��Ͻ]�ϽO�Ͻ��Ͻ��Ͻ��Ͻk�Ͻ��Ͻz�Ͻ��Ͻ��ϽP   P   T�ϽK�Ͻ�Ͻ��Ͻi�Ͻ��Ͻ��Ͻ5�Ͻ��Ͻ_�Ͻ��Ͻ+�Ͻv�ϽZ�Ͻ��Ͻn�Ͻ"�Ͻ�Ͻq�Ͻn�ϽP   P   ��Ͻ��Ͻ��Ͻv�Ͻ��ϽT�ϽU�Ͻ��Ͻ'�Ͻ_�Ͻ��ϽN�Ͻ��Ͻ��Ͻ��Ͻ;�Ͻ��Ͻ7�Ͻ��Ͻ_�ϽP   P   o�Ͻ��Ͻ��Ͻ�Ͻd�Ͻ��ϽT�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ_�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ+�Ͻ��Ͻ��Ͻ�ϽP   P   ��Ͻ��Ͻ|�Ͻ\�Ͻ��Ͻd�Ͻ��Ͻi�Ͻ��ϽJ�Ͻ��Ͻw�Ͻ��ϽD�Ͻa�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻu�Ͻ��Ͻ\�Ͻ�Ͻv�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻs�Ͻ�Ͻ��Ͻ��Ͻ��Ͻd�ϽX�ϽP   P   ��Ͻ��Ͻ��Ͻu�Ͻ|�Ͻ��Ͻ��Ͻ�Ͻd�Ͻ��ϽO�Ͻ��Ͻ��Ͻ��Ͻ[�Ͻ^�Ͻ��Ͻ��Ͻq�Ͻ��ϽP   P   d�Ͻ>�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽK�Ͻq�Ͻ��Ͻ��Ͻc�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽT�Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻ��Ͻ��Ͻv�Ͻ��Ͻ>�Ͻ��Ͻv�Ͻc�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽG�Ͻ��ϽP   P   ��Ͻ��Ͻr�ϽC�Ͻd�Ͻk�Ͻ��Ͻ��Ͻ8�Ͻh�Ͻ��Ͻ�ϽB�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻv�Ͻp�ϽP   P   G�Ͻ�ϽQ�Ͻ{�Ͻ{�Ͻf�Ͻ��Ͻp�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ|�Ͻ.�Ͻn�Ͻ��ϽP�ϽC�Ͻv�ϽP   P   ��Ͻ@�Ͻ6�Ͻj�Ͻo�Ͻ,�Ͻ$�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ^�ϽJ�Ͻ��Ͻ��Ͻ��Ͻ+�Ͻ�ϽP�Ͻ��ϽP   P   ��Ͻ^�Ͻ��Ͻi�Ͻ��Ͻ��Ͻ��ϽE�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻh�Ͻ+�Ͻ��Ͻ��ϽP   P   ��Ͻd�Ͻ��Ͻ��ϽF�Ͻ��Ͻ��Ͻk�Ͻ��Ͻ��Ͻh�Ͻl�Ͻ��Ͻ��Ͻ��ϽU�Ͻ��Ͻ��Ͻn�Ͻ��ϽP   P   ��Ͻ�Ͻ��Ͻ.�Ͻ��ϽE�Ͻ��Ͻ��Ͻh�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ.�Ͻ��ϽP   P   ��Ͻy�Ͻ]�ϽO�ϽJ�ϽG�Ͻb�Ͻ'�Ͻi�ϽW�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ|�Ͻ��ϽP   P   ��Ͻ	�ϽK�Ͻp�ϽV�Ͻ��ϽV�Ͻ��Ͻ��Ͻ|�Ͻ��Ͻd�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽJ�Ͻ��ϽB�ϽP   P   ��Ͻ��Ͻw�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ{�Ͻd�Ͻ��Ͻ��Ͻl�Ͻ��Ͻ^�Ͻ��Ͻ�ϽP   P   c�Ͻ��Ͻ��Ͻ��Ͻ@�Ͻ��Ͻo�Ͻ��Ͻ��Ͻ�Ͻ/�Ͻ�Ͻ��Ͻ��Ͻ��Ͻh�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   v�Ͻ&�Ͻ��Ͻ��ϽE�Ͻ��Ͻ��Ͻx�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ|�ϽW�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻh�ϽP   P   ��Ͻ��Ͻ��ϽZ�ϽV�Ͻ��Ͻ��Ͻ��Ͻ5�Ͻ��Ͻ��Ͻ��Ͻ��Ͻi�Ͻh�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ8�ϽP   P   >�Ͻ��Ͻ��Ͻ��Ͻj�Ͻ��Ͻ{�Ͻ��Ͻ��Ͻx�Ͻ��Ͻ��Ͻ��Ͻ'�Ͻ��Ͻk�ϽE�Ͻ��Ͻp�Ͻ��ϽP   P   ��ϽG�Ͻ��Ͻ��Ͻ|�Ͻu�Ͻ#�Ͻ{�Ͻ��Ͻ��Ͻo�Ͻ��ϽV�Ͻb�Ͻ��Ͻ��Ͻ��Ͻ$�Ͻ��Ͻ��ϽP   P   v�Ͻ%�ϽK�Ͻ��Ͻ��Ͻ	�Ͻu�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽG�ϽE�Ͻ��Ͻ��Ͻ,�Ͻf�Ͻk�ϽP   P   ��ϽP�Ͻ��Ͻ/�Ͻ��Ͻ��Ͻ|�Ͻj�ϽV�ϽE�Ͻ@�Ͻ��ϽV�ϽJ�Ͻ��ϽF�Ͻ��Ͻo�Ͻ{�Ͻd�ϽP   P   ��Ͻ�Ͻ��Ͻ �Ͻ/�Ͻ��Ͻ��Ͻ��ϽZ�Ͻ��Ͻ��Ͻ��Ͻp�ϽO�Ͻ.�Ͻ��Ͻi�Ͻj�Ͻ{�ϽC�ϽP   P   ��Ͻ=�ϽD�Ͻ��Ͻ��ϽK�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻw�ϽK�Ͻ]�Ͻ��Ͻ��Ͻ��Ͻ6�ϽQ�Ͻr�ϽP   P   ��Ͻ��Ͻ=�Ͻ�ϽP�Ͻ%�ϽG�Ͻ��Ͻ��Ͻ&�Ͻ��Ͻ��Ͻ	�Ͻy�Ͻ�Ͻd�Ͻ^�Ͻ@�Ͻ�Ͻ��ϽP   P   ��Ͻ*�ϽL�Ͻe�Ͻ\�Ͻ��Ͻ@�Ͻ*�Ͻ9�Ͻ��Ͻ��Ͻ��Ͻ!�Ͻ�Ͻ3�Ͻ��Ͻ(�Ͻf�Ͻ=�Ͻ-�ϽP   P   -�Ͻ��Ͻ*�Ͻ��Ͻ�Ͻg�ϽD�Ͻ.�Ͻg�Ͻ��Ͻ?�Ͻl�Ͻ��Ͻ��Ͻ7�Ͻ5�Ͻ��Ͻ�Ͻ��Ͻ
�ϽP   P   =�Ͻ7�ϽQ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽL�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   f�Ͻ��Ͻ��Ͻ=�Ͻ%�Ͻ��Ͻ��Ͻ��Ͻ�ϽV�Ͻ��Ͻ��Ͻ��Ͻ��ϽK�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   (�Ͻ��Ͻ�Ͻ��Ͻ.�Ͻ��Ͻ��Ͻ��Ͻ��Ͻx�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��ϽL�ϽO�Ͻ�ϽV�Ͻ��Ͻ9�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ5�ϽP   P   3�Ͻ��ϽD�Ͻ�ϽK�Ͻ��Ͻ,�ϽE�Ͻ��Ͻz�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽK�Ͻ��Ͻ7�ϽP   P   �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   !�Ͻ�Ͻn�ϽO�ϽX�ϽG�Ͻ{�Ͻ �Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ�Ͻl�ϽD�Ͻr�Ͻt�Ͻ3�Ͻm�Ͻ|�Ͻ��Ͻ`�Ͻ:�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽL�Ͻl�ϽP   P   ��Ͻ��Ͻx�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ �Ͻs�Ͻ��Ͻ��Ͻ`�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ?�ϽP   P   ��Ͻ��ϽV�Ͻ:�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ@�Ͻ+�Ͻ��Ͻ��Ͻ��Ͻ��Ͻz�Ͻ��Ͻx�ϽV�Ͻ��Ͻ��ϽP   P   9�ϽZ�Ͻ|�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ~�Ͻ@�Ͻs�Ͻ|�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻg�ϽP   P   *�Ͻ�Ͻ��Ͻ'�Ͻ��Ͻ��Ͻp�Ͻ��Ͻ�Ͻ��Ͻ �Ͻm�Ͻ �Ͻ�ϽE�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ.�ϽP   P   @�ϽV�Ͻ��Ͻ�ϽF�Ͻn�Ͻ�Ͻp�Ͻ��Ͻ��Ͻ�Ͻ3�Ͻ{�Ͻ��Ͻ,�Ͻ9�Ͻ��Ͻ��Ͻ��ϽD�ϽP   P   ��Ͻ��Ͻ��ϽY�ϽT�Ͻ��Ͻn�Ͻ��Ͻ��Ͻ��Ͻ��Ͻt�ϽG�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻg�ϽP   P   \�Ͻ[�ϽZ�Ͻ��Ͻ��ϽT�ϽF�Ͻ��Ͻ��Ͻ��Ͻ�Ͻr�ϽX�Ͻ��ϽK�ϽV�Ͻ.�Ͻ%�Ͻ��Ͻ�ϽP   P   e�Ͻo�Ͻ5�Ͻ0�Ͻ��ϽY�Ͻ�Ͻ'�Ͻ�Ͻ:�Ͻ�ϽD�ϽO�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ=�Ͻ��Ͻ��ϽP   P   L�Ͻ��ϽL�Ͻ5�ϽZ�Ͻ��Ͻ��Ͻ��Ͻ|�ϽV�Ͻx�Ͻl�Ͻn�Ͻ��ϽD�ϽO�Ͻ�Ͻ��ϽQ�Ͻ*�ϽP   P   *�Ͻ��Ͻ��Ͻo�Ͻ[�Ͻ��ϽV�Ͻ�ϽZ�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��ϽL�Ͻ��Ͻ��Ͻ7�Ͻ��ϽP   P   g�ϽK�Ͻ��Ͻm�Ͻu�Ͻ[�Ͻ��Ͻ��Ͻ��ϽT�Ͻ+�ϽG�Ͻ��Ͻ��Ͻ��ϽX�Ͻ��Ͻv�Ͻ��ϽK�ϽP   P   K�ϽE�Ͻ`�Ͻ#�Ͻ��ϽY�Ͻh�Ͻ��Ͻ��Ͻ��ϽS�Ͻ[�Ͻ~�Ͻ��Ͻ��ϽX�ϽO�Ͻd�Ͻ�Ͻr�ϽP   P   ��Ͻ8�Ͻ��Ͻ�Ͻ��Ͻ@�Ͻ�Ͻ&�Ͻ[�Ͻm�Ͻs�Ͻ��Ͻb�Ͻu�Ͻy�ϽH�Ͻ�Ͻ1�Ͻ�Ͻ�ϽP   P   v�Ͻ��Ͻ��ϽW�Ͻ|�ϽM�Ͻc�Ͻ��Ͻ6�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ~�Ͻ��Ͻ!�Ͻ��Ͻi�Ͻ1�Ͻd�ϽP   P   ��Ͻ�Ͻ��Ͻ%�Ͻ��ϽC�Ͻ�Ͻ��Ͻ@�Ͻp�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻc�Ͻ��Ͻ�ϽO�ϽP   P   X�Ͻ��Ͻ��Ͻf�Ͻ��ϽU�ϽP�ϽR�Ͻ!�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ!�ϽH�ϽX�ϽP   P   ��Ͻq�Ͻ(�Ͻ��Ͻ5�ϽV�Ͻ��Ͻ��Ͻv�Ͻ��Ͻ��Ͻv�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻy�Ͻ��ϽP   P   ��Ͻ��Ͻ�ϽH�Ͻp�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻv�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ~�Ͻu�Ͻ��ϽP   P   ��Ͻ��Ͻo�Ͻ4�Ͻ3�Ͻ�Ͻ��Ͻ~�Ͻ��Ͻr�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻb�Ͻ~�ϽP   P   G�Ͻ"�Ͻ��Ͻz�Ͻ@�Ͻb�Ͻ��Ͻc�Ͻ*�Ͻ �ϽT�Ͻ��Ͻ��Ͻ��Ͻv�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ[�ϽP   P   +�ϽP�ϽX�Ͻ��Ͻo�Ͻw�ϽN�Ͻ��Ͻx�ϽC�Ͻa�ϽT�Ͻ��Ͻv�Ͻ��Ͻ��Ͻ��Ͻ��Ͻs�ϽS�ϽP   P   T�ϽC�Ͻ��Ͻw�Ͻy�Ͻ�Ͻ'�Ͻ��Ͻ��Ͻx�ϽC�Ͻ �Ͻr�Ͻ��Ͻ��Ͻ��Ͻp�Ͻ��Ͻm�Ͻ��ϽP   P   ��Ͻ)�Ͻ?�Ͻ��Ͻl�Ͻn�Ͻ/�Ͻe�ϽI�Ͻ��Ͻx�Ͻ*�Ͻ��Ͻ��Ͻv�Ͻ!�Ͻ@�Ͻ6�Ͻ[�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻt�ϽP�Ͻ��ϽX�Ͻe�Ͻ��Ͻ��Ͻc�Ͻ~�Ͻ��Ͻ��ϽR�Ͻ��Ͻ��Ͻ&�Ͻ��ϽP   P   ��Ͻ��ϽK�Ͻ��ϽT�Ͻ<�Ͻ'�Ͻ��Ͻ/�Ͻ'�ϽN�Ͻ��Ͻ��Ͻ��Ͻ��ϽP�Ͻ�Ͻc�Ͻ�Ͻh�ϽP   P   [�Ͻv�Ͻ&�Ͻ;�Ͻc�ϽZ�Ͻ<�ϽP�Ͻn�Ͻ�Ͻw�Ͻb�Ͻ�Ͻ�ϽV�ϽU�ϽC�ϽM�Ͻ@�ϽY�ϽP   P   u�Ͻ��Ͻ��Ͻ]�Ͻ�Ͻc�ϽT�Ͻt�Ͻl�Ͻy�Ͻo�Ͻ@�Ͻ3�Ͻp�Ͻ5�Ͻ��Ͻ��Ͻ|�Ͻ��Ͻ��ϽP   P   m�Ͻ9�Ͻb�Ͻ%�Ͻ]�Ͻ;�Ͻ��Ͻ��Ͻ��Ͻw�Ͻ��Ͻz�Ͻ4�ϽH�Ͻ��Ͻf�Ͻ%�ϽW�Ͻ�Ͻ#�ϽP   P   ��Ͻ��Ͻ��Ͻb�Ͻ��Ͻ&�ϽK�Ͻ��Ͻ?�Ͻ��ϽX�Ͻ��Ͻo�Ͻ�Ͻ(�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ`�ϽP   P   K�ϽW�Ͻ��Ͻ9�Ͻ��Ͻv�Ͻ��Ͻ��Ͻ)�ϽC�ϽP�Ͻ"�Ͻ��Ͻ��Ͻq�Ͻ��Ͻ�Ͻ��Ͻ8�ϽE�ϽP   P   ��Ͻ�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ
�Ͻ��ϽA�Ͻ��Ͻ��Ͻ~�Ͻ{�Ͻ�Ͻ>�Ͻ��ϽR�Ͻ�Ͻ&�Ͻ�ϽP   P   �ϽH�Ͻ,�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ!�ϽF�Ͻ��Ͻ��Ͻs�Ͻ��ϽY�Ͻ��Ͻf�Ͻt�Ͻ��ϽJ�ϽP   P   &�Ͻ7�Ͻ$�Ͻ��Ͻ��Ͻ7�Ͻo�Ͻ��ϽM�Ͻ{�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽE�Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻ/�Ͻ��Ͻi�ϽV�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ<�Ͻ��Ͻ�Ͻk�Ͻl�Ͻ^�ϽE�Ͻt�ϽP   P   R�Ͻ��ϽA�Ͻ��Ͻ)�ϽI�Ͻ��ϽV�Ͻ��Ͻ��Ͻ`�Ͻ��Ͻ��Ͻ��Ͻw�Ͻ��Ͻ��Ͻl�Ͻ��Ͻf�ϽP   P   ��Ͻ��Ͻ}�Ͻx�Ͻ �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻk�Ͻ��Ͻ��ϽP   P   >�Ͻ�Ͻ��Ͻ{�Ͻ��Ͻ��Ͻc�Ͻ[�Ͻ{�Ͻ��Ͻu�Ͻ��Ͻ��Ͻ��Ͻ'�Ͻ��Ͻw�Ͻ�Ͻ��ϽY�ϽP   P   �Ͻ��Ͻ �ϽL�Ͻi�ϽC�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   {�Ͻ_�Ͻ2�Ͻ��ϽQ�ϽK�Ͻ2�ϽN�Ͻ��Ͻ?�Ͻ��Ͻ'�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ<�Ͻ��Ͻs�ϽP   P   ~�Ͻ�Ͻ�Ͻ
�Ͻ�Ͻ9�ϽF�Ͻ��Ͻ��Ͻp�Ͻ��Ͻ��Ͻ'�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ4�Ͻ,�Ͻ*�Ͻ�Ͻ�Ͻ�Ͻ_�ϽC�Ͻ��Ͻ��Ͻ��Ͻ��Ͻu�Ͻ�Ͻ`�Ͻ��Ͻ��Ͻ��ϽP   P   ��ϽB�Ͻ?�Ͻ��Ͻ��Ͻ��Ͻ+�Ͻ��Ͻ�Ͻ.�ϽC�Ͻp�Ͻ?�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ{�ϽF�ϽP   P   A�Ͻ��Ͻ2�Ͻ:�Ͻ~�Ͻx�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ_�Ͻ��Ͻ��Ͻ��Ͻ{�Ͻ��Ͻ��Ͻ��ϽM�Ͻ!�ϽP   P   ��Ͻ}�Ͻ&�Ͻ�Ͻ��Ͻ]�Ͻ��Ͻw�Ͻ��Ͻ��Ͻ�Ͻ��ϽN�Ͻ��Ͻ[�Ͻ��ϽV�Ͻ��Ͻ��Ͻ��ϽP   P   
�Ͻ>�Ͻ��ϽR�Ͻ��ϽZ�Ͻt�Ͻ��Ͻ��Ͻ+�Ͻ�ϽF�Ͻ2�Ͻ�Ͻc�Ͻ��Ͻ��ϽV�Ͻo�Ͻ��ϽP   P   ��Ͻ�ϽE�Ͻ��ϽV�Ͻ��ϽZ�Ͻ]�Ͻx�Ͻ��Ͻ�Ͻ9�ϽK�ϽC�Ͻ��Ͻ��ϽI�Ͻi�Ͻ7�Ͻ��ϽP   P   ��Ͻ.�ϽK�Ͻu�Ͻ��ϽV�Ͻ��Ͻ��Ͻ~�Ͻ��Ͻ*�Ͻ�ϽQ�Ͻi�Ͻ��Ͻ �Ͻ)�Ͻ��Ͻ��Ͻ��ϽP   P   �Ͻ@�Ͻ��Ͻ��Ͻu�Ͻ��ϽR�Ͻ�Ͻ:�Ͻ��Ͻ,�Ͻ
�Ͻ��ϽL�Ͻ{�Ͻx�Ͻ��Ͻ/�Ͻ��Ͻ�ϽP   P   �Ͻz�Ͻ�Ͻ��ϽK�ϽE�Ͻ��Ͻ&�Ͻ2�Ͻ?�Ͻ4�Ͻ�Ͻ2�Ͻ �Ͻ��Ͻ}�ϽA�Ͻ��Ͻ$�Ͻ,�ϽP   P   �Ͻv�Ͻz�Ͻ@�Ͻ.�Ͻ�Ͻ>�Ͻ}�Ͻ��ϽB�Ͻ��Ͻ�Ͻ_�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ7�ϽH�ϽP   P   &�Ͻ�Ͻ��Ͻ�Ͻ,�Ͻ��Ͻ<�Ͻ_�Ͻ�Ͻ?�Ͻ-�Ͻ�ϽH�Ͻ��Ͻ_�Ͻ]�Ͻ��Ͻ
�Ͻ��Ͻ�ϽP   P   �Ͻ3�Ͻ6�Ͻv�Ͻ��Ͻ�Ͻ��ϽL�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ0�Ͻ��Ͻ�Ͻ��Ͻc�Ͻ6�ϽP   P   ��Ͻ�Ͻ��Ͻn�Ͻ�Ͻ�Ͻ2�Ͻ4�Ͻ}�Ͻ��Ͻ��Ͻ7�Ͻ��Ͻ��Ͻ��Ͻ6�ϽN�Ͻ�Ͻ]�Ͻc�ϽP   P   
�Ͻ�Ͻ5�Ͻ-�Ͻ��Ͻ�Ͻ��ϽQ�Ͻy�Ͻ?�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ#�Ͻj�Ͻ7�Ͻ��Ͻ�Ͻ��ϽP   P   ��ϽA�Ͻ@�Ͻ.�Ͻ-�Ͻ�Ͻ?�Ͻ8�ϽH�Ͻz�Ͻf�Ͻ��Ͻ�Ͻ��Ͻ��Ͻi�Ͻ}�Ͻ7�ϽN�Ͻ�ϽP   P   ]�Ͻ�Ͻ��Ͻ��Ͻb�Ͻ��Ͻ��Ͻ:�Ͻ��Ͻ��Ͻ(�Ͻ�Ͻ��Ͻd�Ͻ��Ͻ3�Ͻi�Ͻj�Ͻ6�Ͻ��ϽP   P   _�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��ϽE�ϽG�Ͻ��Ͻ!�Ͻ��Ͻ��Ͻ`�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ#�Ͻ��Ͻ0�ϽP   P   ��Ͻy�Ͻ+�Ͻ��Ͻ��Ͻ\�Ͻ��Ͻ}�Ͻ��Ͻ��Ͻ��Ͻ��Ͻq�Ͻ��Ͻ��Ͻd�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   H�Ͻ�Ͻa�Ͻ9�Ͻ��Ͻ�ϽE�Ͻ�Ͻ7�Ͻ��Ͻ��Ͻ(�Ͻ��Ͻq�Ͻ`�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��ϽP   P   �Ͻ+�ϽC�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ0�ϽE�Ͻ�Ͻ��Ͻ6�Ͻ(�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ7�Ͻ��ϽP   P   -�Ͻj�ϽC�Ͻ)�Ͻ��Ͻ��ϽU�Ͻ7�Ͻ>�ϽW�Ͻ6�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ(�Ͻf�Ͻ��Ͻ��Ͻ��ϽP   P   ?�ϽK�Ͻ �Ͻ{�Ͻ��Ͻ��Ͻ��Ͻi�Ͻ�Ͻ�ϽW�Ͻ�Ͻ��Ͻ��Ͻ!�Ͻ��Ͻz�Ͻ?�Ͻ��Ͻ��ϽP   P   �Ͻ0�ϽB�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ>�ϽE�Ͻ7�Ͻ��Ͻ��Ͻ��ϽH�Ͻy�Ͻ}�Ͻ�ϽP   P   _�ϽN�Ͻ;�Ͻ!�Ͻq�Ͻ��Ͻ�Ͻ��Ͻ��Ͻi�Ͻ7�Ͻ0�Ͻ�Ͻ}�ϽG�Ͻ:�Ͻ8�ϽQ�Ͻ4�ϽL�ϽP   P   <�Ͻ��Ͻ�Ͻ��ϽU�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��ϽU�Ͻ��ϽE�Ͻ��ϽE�Ͻ��Ͻ?�Ͻ��Ͻ2�Ͻ��ϽP   P   ��Ͻ��ϽL�ϽK�Ͻ �ϽV�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ\�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�Ͻ�ϽP   P   ,�ϽA�Ͻ��Ͻ��Ͻ��Ͻ �ϽU�Ͻq�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻb�Ͻ-�Ͻ��Ͻ�Ͻ��ϽP   P   �Ͻh�Ͻ��Ͻ��Ͻ��ϽK�Ͻ��Ͻ!�Ͻ��Ͻ{�Ͻ)�Ͻ��Ͻ9�Ͻ��Ͻ��Ͻ��Ͻ.�Ͻ-�Ͻn�Ͻv�ϽP   P   ��Ͻ,�Ͻ�Ͻ��Ͻ��ϽL�Ͻ�Ͻ;�ϽB�Ͻ �ϽC�ϽC�Ͻa�Ͻ+�Ͻ�Ͻ��Ͻ@�Ͻ5�Ͻ��Ͻ6�ϽP   P   �Ͻ��Ͻ,�Ͻh�ϽA�Ͻ��Ͻ��ϽN�Ͻ0�ϽK�Ͻj�Ͻ+�Ͻ�Ͻy�Ͻ��Ͻ�ϽA�Ͻ�Ͻ�Ͻ3�ϽP   P   ?�Ͻ�Ͻ�Ͻ �Ͻ�Ͻ1�Ͻ5�ϽL�Ͻ<�Ͻ��Ͻ��Ͻ��ϽJ�Ͻb�Ͻ	�Ͻ�Ͻ	�Ͻ�Ͻ6�Ͻ�ϽP   P   �Ͻ�Ͻ��Ͻ��Ͻ��Ͻb�Ͻ*�Ͻ]�ϽQ�Ͻ|�Ͻ��Ͻ	�ϽV�ϽT�ϽK�ϽF�Ͻ|�Ͻ��Ͻ��Ͻ@�ϽP   P   6�Ͻn�Ͻ��Ͻ��Ͻ��Ͻb�Ͻ]�Ͻ��Ͻn�Ͻ��Ͻ{�Ͻ��Ͻ��Ͻ �Ͻn�Ͻ~�ϽQ�ϽT�Ͻ��Ͻ��ϽP   P   �ϽY�Ͻ��Ͻ'�Ͻ��ϽJ�Ͻ�Ͻj�Ͻ��Ͻ��Ͻ��Ͻ��Ͻe�Ͻ��Ͻ��Ͻ��Ͻk�Ͻ�ϽT�Ͻ��ϽP   P   	�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽE�Ͻ��Ͻ��Ͻ��Ͻ�Ͻm�Ͻ��Ͻr�Ͻ�Ͻ��Ͻ��Ͻk�ϽQ�Ͻ|�ϽP   P   �Ͻ��Ͻj�ϽP�Ͻ��Ͻ'�ϽG�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻl�Ͻk�Ͻ|�Ͻ��Ͻ��Ͻ��Ͻ~�ϽF�ϽP   P   	�Ͻ��Ͻ)�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ=�Ͻ��Ͻ��Ͻ��Ͻ��ϽY�Ͻ�Ͻ|�Ͻ�Ͻ��Ͻn�ϽK�ϽP   P   b�Ͻ��Ͻ��ϽT�ϽU�Ͻ��Ͻ��Ͻg�Ͻ[�Ͻ��Ͻ��Ͻp�Ͻo�Ͻ��ϽY�Ͻk�Ͻr�Ͻ��Ͻ �ϽT�ϽP   P   J�Ͻ��Ͻ�Ͻ��Ͻ]�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��ϽP�Ͻ��Ͻ��Ͻo�Ͻ��Ͻl�Ͻ��Ͻe�Ͻ��ϽV�ϽP   P   ��Ͻ&�Ͻw�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ7�Ͻ��Ͻ�Ͻ��Ͻ��Ͻp�Ͻ��Ͻ��Ͻm�Ͻ��Ͻ��Ͻ	�ϽP   P   ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽC�Ͻr�Ͻ�ϽP�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ{�Ͻ��ϽP   P   ��ϽK�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽC�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ|�ϽP   P   <�Ͻ��Ͻ �Ͻg�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ7�Ͻ�Ͻ[�Ͻ=�Ͻ��Ͻ��Ͻ��Ͻn�ϽQ�ϽP   P   L�Ͻ0�Ͻg�Ͻ��Ͻ��Ͻ��Ͻ`�Ͻe�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻg�Ͻ��Ͻ��Ͻ��Ͻj�Ͻ��Ͻ]�ϽP   P   5�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ`�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��ϽG�ϽE�Ͻ�Ͻ]�Ͻ*�ϽP   P   1�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ'�Ͻ��ϽJ�Ͻb�Ͻb�ϽP   P   �Ͻ��ϽW�ϽR�Ͻ[�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ]�ϽU�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P    �Ͻ��Ͻt�Ͻ��ϽR�Ͻ�Ͻ��Ͻ��Ͻg�Ͻ��Ͻ��Ͻ�Ͻ��ϽT�Ͻ��ϽP�Ͻ��Ͻ'�Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻt�ϽW�Ͻ��Ͻ�Ͻg�Ͻ �Ͻ�Ͻ�Ͻw�Ͻ�Ͻ��Ͻ)�Ͻj�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   �Ͻ^�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ0�Ͻ��ϽK�Ͻ�Ͻ&�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽY�Ͻn�Ͻ�ϽP   P   }�Ͻ~�Ͻ��Ͻ��Ͻ��Ͻ��Ͻb�Ͻ��Ͻ��Ͻ/�Ͻ��Ͻ^�ϽL�Ͻ��Ͻ�Ͻ��Ͻp�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻj�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ0�Ͻ�Ͻ�Ͻo�ϽD�Ͻ:�ϽG�ϽD�ϽG�ϽW�Ͻ��Ͻ�Ͻ��Ͻu�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�Ͻ]�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ-�ϽP�ϽO�Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ �Ͻ��Ͻ��ϽS�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ
�Ͻ��Ͻ��ϽI�Ͻo�Ͻ��Ͻ�Ͻ�ϽP   P   p�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ/�Ͻ#�Ͻ$�Ͻ��Ͻ��Ͻ|�Ͻo�Ͻ��Ͻ��ϽP   P   ��Ͻ �ϽX�Ͻj�Ͻ��Ͻ��ϽM�Ͻ?�Ͻ"�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ(�Ͻ:�Ͻ��Ͻ��ϽI�ϽO�ϽW�ϽP   P   �ϽF�Ͻ��Ͻ��Ͻ��ϽS�Ͻ �ϽC�Ͻf�Ͻ�Ͻ��ϽA�Ͻ�Ͻm�Ͻ�Ͻ:�Ͻ��Ͻ��ϽP�ϽG�ϽP   P   ��ϽW�ϽZ�Ͻg�Ͻ5�Ͻ]�ϽU�Ͻ��Ͻ7�Ͻ
�Ͻ�Ͻ!�Ͻ�ϽY�Ͻm�Ͻ(�Ͻ$�Ͻ��Ͻ-�ϽD�ϽP   P   L�Ͻ �Ͻ��Ͻ��Ͻs�Ͻ��Ͻ��Ͻ!�ϽD�Ͻy�Ͻ��Ͻ�Ͻ%�Ͻ�Ͻ�Ͻ�Ͻ#�Ͻ
�Ͻ��ϽG�ϽP   P   ^�Ͻ �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ'�ϽC�Ͻ@�Ͻ��Ͻ�Ͻ!�ϽA�Ͻ�Ͻ/�Ͻ�Ͻ��Ͻ:�ϽP   P   ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ
�Ͻ��Ͻ�Ͻ��Ͻ@�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽD�ϽP   P   /�Ͻ�Ͻ��Ͻ7�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ2�Ͻ��Ͻ�ϽC�Ͻy�Ͻ
�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻo�ϽP   P   ��Ͻ�Ͻ�Ͻ�Ͻ
�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ2�Ͻ��Ͻ'�ϽD�Ͻ7�Ͻf�Ͻ"�Ͻ��Ͻ�Ͻ��Ͻ�ϽP   P   ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ
�Ͻ��Ͻ!�Ͻ��ϽC�Ͻ?�Ͻ��ϽS�Ͻ]�Ͻ�ϽP   P   b�Ͻ'�Ͻ!�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽU�Ͻ �ϽM�Ͻ��Ͻ��Ͻ�Ͻ0�ϽP   P   ��Ͻ$�Ͻ@�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ]�ϽS�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ��Ͻ�ϽA�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ
�Ͻ��Ͻ��Ͻ��Ͻs�Ͻ5�Ͻ��Ͻ��Ͻ��Ͻ �Ͻ�Ͻ��ϽP   P   ��Ͻ��Ͻj�Ͻ��ϽA�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ7�Ͻ��Ͻ��Ͻ��Ͻg�Ͻ��Ͻj�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ4�Ͻj�Ͻ�Ͻ@�Ͻ!�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��ϽZ�Ͻ��ϽX�Ͻ�Ͻ��Ͻ��Ͻ��ϽP   P   ~�Ͻx�Ͻ��Ͻ��Ͻ��Ͻ$�Ͻ'�Ͻ�Ͻ�Ͻ�Ͻ��Ͻ �Ͻ �ϽW�ϽF�Ͻ �Ͻ��Ͻ��Ͻ��Ͻj�ϽP   P   2�Ͻp�ϽX�ϽC�Ͻ�Ͻ��Ͻ�Ͻ<�Ͻa�Ͻ/�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ6�ϽJ�Ͻn�ϽP   P   n�Ͻg�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ2�Ͻ��ϽZ�Ͻ��Ͻ}�Ͻz�Ͻ��Ͻe�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   J�Ͻ��Ͻ�Ͻm�Ͻv�Ͻ��ϽP�Ͻ`�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻd�Ͻd�Ͻ�Ͻ��Ͻ�Ͻ��ϽP   P   6�Ͻ��Ͻu�Ͻ3�Ͻ��Ͻ��Ͻ|�Ͻd�Ͻz�ϽA�Ͻ_�Ͻ��Ͻ;�Ͻ4�Ͻh�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻg�Ͻx�Ͻ�Ͻ��ϽW�Ͻ��Ͻ��ϽN�Ͻ��Ͻl�Ͻ�ϽI�Ͻ��Ͻk�Ͻn�Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ&�Ͻx�Ͻ��Ͻ��Ͻ��Ͻ	�ϽW�Ͻ]�Ͻ>�Ͻh�ϽT�Ͻ��Ͻ��Ͻ��Ͻ0�Ͻk�Ͻ��Ͻd�Ͻ��ϽP   P   ��Ͻ`�Ͻ��ϽT�Ͻ��Ͻh�Ͻ��Ͻ*�Ͻ��Ͻe�Ͻ��Ͻy�Ͻ��Ͻk�Ͻ��Ͻ��Ͻ��Ͻh�Ͻd�Ͻe�ϽP   P   �Ͻ��Ͻ��Ͻ:�Ͻ��Ͻ��Ͻ��Ͻ#�Ͻ��Ͻ��ϽN�Ͻ@�Ͻ��Ͻ7�Ͻk�Ͻ��ϽI�Ͻ4�Ͻ��Ͻ��ϽP   P   �Ͻ9�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽZ�Ͻm�Ͻ��Ͻ�Ͻ<�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ;�Ͻ��Ͻz�ϽP   P   ��Ͻ,�Ͻ��Ͻ��Ͻ��Ͻ��Ͻp�Ͻ��Ͻ
�ϽY�Ͻ��Ͻ��Ͻ�Ͻ@�Ͻy�ϽT�Ͻl�Ͻ��Ͻ��Ͻ}�ϽP   P   ��Ͻ,�Ͻ��Ͻ��ϽG�Ͻv�Ͻu�Ͻ��Ͻ��Ͻ&�Ͻ��Ͻ��Ͻ��ϽN�Ͻ��Ͻh�Ͻ��Ͻ_�Ͻ��Ͻ��ϽP   P   /�Ͻ7�ϽY�Ͻ_�Ͻ-�Ͻ.�Ͻ�ϽK�ϽU�ϽW�Ͻ&�ϽY�Ͻm�Ͻ��Ͻe�Ͻ>�ϽN�ϽA�Ͻ��ϽZ�ϽP   P   a�ϽM�Ͻ��Ͻ\�ϽE�Ͻ^�Ͻf�ϽI�ϽK�ϽU�Ͻ��Ͻ
�ϽZ�Ͻ��Ͻ��Ͻ]�Ͻ��Ͻz�Ͻ��Ͻ��ϽP   P   <�Ͻ��Ͻ��Ͻ��ϽU�ϽE�Ͻ2�Ͻ[�ϽI�ϽK�Ͻ��Ͻ��Ͻ�Ͻ#�Ͻ*�ϽW�Ͻ��Ͻd�Ͻ`�Ͻ2�ϽP   P   �Ͻ��Ͻ��Ͻ��ϽN�Ͻ�Ͻ��Ͻ2�Ͻf�Ͻ�Ͻu�Ͻp�Ͻ��Ͻ��Ͻ��Ͻ	�ϽW�Ͻ|�ϽP�Ͻ��ϽP   P   ��Ͻ_�Ͻ��Ͻh�Ͻ��Ͻ��Ͻ�ϽE�Ͻ^�Ͻ.�Ͻv�Ͻ��Ͻ��Ͻ��Ͻh�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽN�ϽU�ϽE�Ͻ-�ϽG�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻv�Ͻ��ϽP   P   C�Ͻi�Ͻ��Ͻ%�Ͻ�Ͻh�Ͻ��Ͻ��Ͻ\�Ͻ_�Ͻ��Ͻ��Ͻ��Ͻ:�ϽT�Ͻ��Ͻx�Ͻ3�Ͻm�Ͻ��ϽP   P   X�Ͻ{�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽY�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻx�Ͻg�Ͻu�Ͻ�Ͻ��ϽP   P   p�Ͻ'�Ͻ{�Ͻi�Ͻ��Ͻ_�Ͻ��Ͻ��ϽM�Ͻ7�Ͻ,�Ͻ,�Ͻ9�Ͻ��Ͻ`�Ͻ&�Ͻ��Ͻ��Ͻ��Ͻg�ϽP   P   ��Ͻ��Ͻ@�ϽY�ϽR�Ͻ��Ͻ��Ͻ'�Ͻ�Ͻ��Ͻ9�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ �ϽE�Ͻ6�Ͻ��ϽP   P   ��Ͻ��Ͻ��ϽK�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ:�Ͻj�Ͻ�Ͻ��Ͻ��ϽH�Ͻ1�Ͻ��Ͻ��Ͻ��Ͻ0�Ͻ��ϽP   P   6�Ͻ��Ͻo�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ]�Ͻ��Ͻ��Ͻ:�Ͻ��ϽH�Ͻ��Ͻd�Ͻb�Ͻ��Ͻ��Ͻa�Ͻ0�ϽP   P   E�Ͻo�Ͻ2�ϽX�Ͻ��Ͻ��Ͻ��Ͻ.�Ͻ8�ϽY�Ͻ��Ͻ�ϽK�Ͻ��Ͻs�Ͻ4�Ͻ8�Ͻ��Ͻ��Ͻ��ϽP   P    �Ͻ�Ͻ��Ͻ#�Ͻn�Ͻ��Ͻ�Ͻ*�Ͻp�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ+�Ͻ8�Ͻ��Ͻ��ϽP   P   ��ϽU�ϽU�Ͻ��Ͻ�Ͻ��Ͻ��ϽF�Ͻ�Ͻ��Ͻ�ϽN�Ͻ�Ͻ
�Ͻ��Ͻ��Ͻ��Ͻ4�Ͻb�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻx�Ͻ�Ͻ��Ͻ$�Ͻ��Ͻ��Ͻd�Ͻ��Ͻe�Ͻa�Ͻ�Ͻ7�Ͻ��Ͻ��Ͻs�Ͻd�Ͻ1�ϽP   P   �Ͻ��Ͻb�Ͻ.�Ͻ��Ͻc�Ͻ��Ͻ(�ϽE�ϽS�Ͻ��Ͻ��Ͻ�ϽZ�Ͻ�Ͻ
�Ͻ��Ͻ��Ͻ��ϽH�ϽP   P   ��Ͻ��Ͻ��Ͻf�Ͻ-�Ͻp�Ͻ��Ͻ��Ͻ �ϽY�Ͻ��Ͻ�Ͻ��Ͻ�Ͻa�Ͻ�Ͻ��ϽK�ϽH�Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻ��Ͻ4�Ͻ%�ϽS�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻe�ϽN�Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   9�Ͻ��Ͻ��Ͻw�Ͻ$�Ͻ|�ϽG�ϽW�Ͻ �Ͻ��ϽR�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ:�Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻz�Ͻ��Ͻ��Ͻp�Ͻ��Ͻ��Ͻ��Ͻ�ϽY�ϽS�Ͻd�Ͻ��Ͻ��ϽY�Ͻ��Ͻj�ϽP   P   �Ͻ�Ͻ��Ͻ��Ͻ��Ͻ �Ͻ��Ͻ�Ͻ��Ͻ��Ͻ �Ͻ��Ͻ �ϽE�Ͻ��Ͻ�Ͻp�Ͻ8�Ͻ��Ͻ:�ϽP   P   '�Ͻ��Ͻ��Ͻc�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻp�ϽW�Ͻ��Ͻ��Ͻ(�Ͻ��ϽF�Ͻ*�Ͻ.�Ͻ]�Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽG�ϽS�Ͻ��Ͻ��Ͻ$�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ��Ͻc�ϽD�Ͻ6�Ͻ��Ͻ��Ͻ�Ͻ �Ͻ��Ͻ|�Ͻ%�Ͻp�Ͻc�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   R�Ͻ;�Ͻ��Ͻ"�ϽF�Ͻ6�Ͻ�Ͻ��Ͻ��Ͻz�Ͻ$�Ͻ4�Ͻ-�Ͻ��Ͻ�Ͻ�Ͻn�Ͻ��Ͻ��Ͻ��ϽP   P   Y�Ͻ#�Ͻx�Ͻ��Ͻ"�ϽD�Ͻ��Ͻc�Ͻ��Ͻ��Ͻw�Ͻ��Ͻf�Ͻ.�Ͻx�Ͻ��Ͻ#�ϽX�Ͻ�ϽK�ϽP   P   @�ϽE�Ͻ��Ͻx�Ͻ��Ͻc�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻb�Ͻ��ϽU�Ͻ��Ͻ2�Ͻo�Ͻ��ϽP   P   ��Ͻ��ϽE�Ͻ#�Ͻ;�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽU�Ͻ�Ͻo�Ͻ��Ͻ��ϽP   P   	�Ͻ�Ͻ��Ͻ�Ͻ��Ͻf�Ͻx�Ͻ��Ͻ��Ͻ��Ͻ#�Ͻz�Ͻ��Ͻ��Ͻ��ϽY�Ͻ �Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ{�Ͻ��Ͻc�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ6�Ͻ��Ͻc�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻd�Ͻ��Ͻ��ϽN�Ͻ��Ͻ��Ͻ3�Ͻ��Ͻ��Ͻ(�Ͻ�Ͻ7�Ͻ��Ͻ��Ͻ-�Ͻ�Ͻ~�Ͻj�Ͻ��ϽP   P   �Ͻl�ϽY�Ͻ��Ͻ!�Ͻ��Ͻ �Ͻ��Ͻ��Ͻ+�Ͻ~�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ~�Ͻ��ϽP   P    �Ͻ`�Ͻ�Ͻz�Ͻ��Ͻ`�Ͻ�Ͻ��ϽO�Ͻ"�Ͻ��Ͻ\�Ͻ��ϽE�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻc�ϽP   P   Y�Ͻ@�Ͻ��Ͻ��Ͻ=�Ͻ\�Ͻ�Ͻ'�Ͻ��Ͻ�Ͻ,�Ͻi�Ͻ��Ͻ��ϽI�Ͻ>�Ͻ�Ͻ��Ͻ-�Ͻ��ϽP   P   ��Ͻ��Ͻj�Ͻg�Ͻ`�Ͻ��Ͻw�Ͻ;�Ͻ��Ͻ�Ͻ��ϽS�Ͻ��Ͻe�Ͻ��ϽI�Ͻ��Ͻ�Ͻ��Ͻ6�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻw�Ͻ��Ͻ��Ͻ��Ͻ��ϽF�Ͻ��Ͻs�Ͻe�Ͻ��ϽE�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ&�Ͻ �ϽP�Ͻ
�Ͻ7�Ͻ��Ͻm�Ͻ��ϽG�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ7�Ͻ��ϽP   P   z�Ͻ��ϽT�Ͻ�Ͻ$�Ͻ�Ͻ2�Ͻ �Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽF�ϽS�Ͻi�Ͻ\�Ͻ��Ͻ�Ͻ��ϽP   P   #�Ͻ��ϽI�Ͻ��Ͻ��ϽU�Ͻ��Ͻ��Ͻg�Ͻ��Ͻ��Ͻ��ϽG�Ͻ��Ͻ��Ͻ,�Ͻ��Ͻ~�Ͻ(�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ"�Ͻ+�Ͻ��Ͻ�ϽP   P   ��Ͻ��ϽF�Ͻ��Ͻx�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻg�Ͻ��Ͻm�Ͻ��Ͻ��Ͻ��ϽO�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ=�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ �Ͻ��Ͻ��Ͻ;�Ͻ'�Ͻ��Ͻ��Ͻ3�Ͻc�ϽP   P   x�Ͻ��Ͻ�Ͻ%�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ2�Ͻ7�Ͻw�Ͻw�Ͻ�Ͻ�Ͻ �Ͻ��Ͻ��ϽP   P   f�Ͻ��Ͻ��Ͻ�Ͻ"�Ͻ[�Ͻ��Ͻ��Ͻ��Ͻ��ϽU�Ͻ�Ͻ
�Ͻ��Ͻ��Ͻ\�Ͻ`�Ͻ��Ͻ��Ͻ{�ϽP   P   ��ϽZ�Ͻ3�Ͻ�Ͻ,�Ͻ"�Ͻ��Ͻ��Ͻx�Ͻ��Ͻ��Ͻ$�ϽP�Ͻ�Ͻ`�Ͻ=�Ͻ��Ͻ!�ϽN�Ͻ�ϽP   P   �Ͻs�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ%�Ͻ��Ͻ��Ͻ �Ͻ��Ͻ�Ͻ �Ͻ��Ͻg�Ͻ��Ͻz�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ{�Ͻ��Ͻ��Ͻ3�Ͻ��Ͻ�Ͻ=�ϽF�Ͻ��ϽI�ϽT�Ͻ&�Ͻ��Ͻj�Ͻ��Ͻ�ϽY�Ͻ��Ͻ��ϽP   P   �ϽZ�Ͻ{�Ͻs�ϽZ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ@�Ͻ`�Ͻl�Ͻd�Ͻ��ϽP   P   B�Ͻ��Ͻ-�Ͻf�Ͻ��Ͻ`�ϽW�Ͻ��Ͻ{�Ͻt�Ͻ��Ͻ)�Ͻ��Ͻ��Ͻ��ϽJ�ϽF�Ͻu�Ͻ<�Ͻ��ϽP   P   ��Ͻ��Ͻo�ϽY�Ͻ��Ͻ��Ͻ��Ͻr�ϽM�Ͻ��Ͻ/ н� н��Ͻ7�Ͻ!�Ͻ��Ͻn�Ͻ��Ͻg�Ͻ:�ϽP   P   <�ϽH�Ͻ=�Ͻ}�Ͻ��Ͻ^�Ͻ��Ͻ��Ͻ9 н� нc н� нo нf н� нs�Ͻ�Ͻl�Ͻ�Ͻg�ϽP   P   u�Ͻm�Ͻ��ϽT�Ͻ��Ͻn�Ͻ3�Ͻm�Ͻ��Ͻ� н� н�нnнKн� н��Ͻ>�Ͻ��Ͻl�Ͻ��ϽP   P   F�Ͻ0�Ͻp�Ͻd�Ͻ��Ͻ��Ͻ��ϽD�Ͻ{ н@нeн�нн�нlнн� н>�Ͻ�Ͻn�ϽP   P   J�ϽP�Ͻ��ϽF�Ͻ��ϽC�Ͻ�Ͻ��Ͻ, н1н�н�н�н�н�н�нн��Ͻs�Ͻ��ϽP   P   ��ϽQ�Ͻ��Ͻ �Ͻ��Ͻw�ϽG�Ͻg�Ͻ	 н� нvн�ннqн'н�нlн� н� н!�ϽP   P   ��Ͻ*�Ͻu�Ͻ��Ͻ�Ͻ>�ϽJ�Ͻ��Ͻs�Ͻ� н н�н�н�нqн�н�нKнf н7�ϽP   P   ��Ͻ��Ͻ%�Ͻf�Ͻ��ϽS�Ͻ�Ͻ�Ͻ`�Ͻ��Ͻ# н�н#н�нн�ннnнo н��ϽP   P   )�Ͻ��Ͻv�Ͻ��Ͻ��Ͻf�Ͻ��Ͻ!�Ͻ��Ͻs�Ͻn н� н�н�н�н�н�н�н� н� нP   P   ��Ͻ��Ͻ4�Ͻ��Ͻ��Ͻ|�Ͻ��Ͻ�Ͻ3�Ͻ��Ͻ��Ͻn н# н нvн�нeн� нc н/ нP   P   t�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ;�Ͻs�Ͻ�Ͻ��Ͻ��Ͻs�Ͻ��Ͻ� н� н1н@н� н� н��ϽP   P   {�Ͻ��ϽB�Ͻ�ϽX�Ͻ�Ͻ?�Ͻ(�Ͻn�Ͻ�Ͻ3�Ͻ��Ͻ`�Ͻs�Ͻ	 н, н{ н��Ͻ9 нM�ϽP   P   ��Ͻ�Ͻf�Ͻ%�Ͻt�ϽC�Ͻ�Ͻ��Ͻ(�Ͻs�Ͻ�Ͻ!�Ͻ�Ͻ��Ͻg�Ͻ��ϽD�Ͻm�Ͻ��Ͻr�ϽP   P   W�Ͻ5�Ͻ��Ͻ��Ͻ��Ͻ,�Ͻ��Ͻ�Ͻ?�Ͻ;�Ͻ��Ͻ��Ͻ�ϽJ�ϽG�Ͻ�Ͻ��Ͻ3�Ͻ��Ͻ��ϽP   P   `�Ͻj�Ͻl�Ͻ��Ͻ��Ͻv�Ͻ,�ϽC�Ͻ�Ͻ�Ͻ|�Ͻf�ϽS�Ͻ>�Ͻw�ϽC�Ͻ��Ͻn�Ͻ^�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��ϽO�Ͻ��Ͻ��Ͻt�ϽX�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   f�Ͻh�Ͻ�ϽM�Ͻ��Ͻ��Ͻ��Ͻ%�Ͻ�Ͻ�Ͻ��Ͻ��Ͻf�Ͻ��Ͻ �ϽF�Ͻd�ϽT�Ͻ}�ϽY�ϽP   P   -�Ͻ��Ͻ@�Ͻ�Ͻ��Ͻl�Ͻ��Ͻf�ϽB�Ͻ��Ͻ4�Ͻv�Ͻ%�Ͻu�Ͻ��Ͻ��Ͻp�Ͻ��Ͻ=�Ͻo�ϽP   P   ��Ͻ�Ͻ��Ͻh�Ͻ��Ͻj�Ͻ5�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ*�ϽQ�ϽP�Ͻ0�Ͻm�ϽH�Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻ��ϽL�Ͻ" н� н;н�нн� н1н�нSн� н н��Ͻ��Ͻ��Ͻ}�ϽP   P   }�Ͻq�Ͻa�Ͻ��Ͻ��Ͻ��ϽM нн�н�ннWн�н�н� н@ н��Ͻr�Ͻ��Ͻe�ϽP   P   ��Ͻ��Ͻ��Ͻ�Ͻ}�Ͻ��Ͻ� н�нн�н8н\нн�н[н�н� н н��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ  н)н�н�нPн�нsнDн�нDнzн�н� н нr�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻq�Ͻ��Ͻ� н�нLнUн*н.н�н4нн<н�н�н� н��ϽP   P    н��ϽR�Ͻ/�Ͻ��Ͻ нH нн�нZн�н"н\нhн�н�н<нzн�н@ нP   P   � н нR�Ͻ��ϽH�Ͻ+ н� нн�н%н0н	нAнeнbн�ннDн[н� нP   P   SнE н��Ͻ��Ͻ��Ͻ��Ͻg н+н�нAн�н3нTн�нeнhн4н�н�н�нP   P   �н н��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ7 нн�н�нeн�нTнAн\н�нDнн�нP   P   1н� н��Ͻ��Ͻ��Ͻ��Ͻ,�Ͻu�Ͻ� нSнEн�нeн3н	н"н.нsн\нWнP   P   � н� н
 н��Ͻ��Ͻ&�Ͻ��Ͻ�Ͻ н� н� нEн�н�н0н�н*н�н8ннP   P   н� н��Ͻ]�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ`�Ͻ��Ͻ� нSн�нAн%нZнUнPн�н�нP   P   �нt н нq�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ`�Ͻ н� нн�н�н�нLн�нн�нP   P   ;нO н��Ͻ��Ͻ��Ͻ��Ͻ6�Ͻ��Ͻ��Ͻ��Ͻ�Ͻu�Ͻ7 н+ннн�н�н�ннP   P   � нl н��Ͻ�Ͻ��Ͻ��Ͻ`�Ͻ6�Ͻ��Ͻ��Ͻ��Ͻ,�Ͻ��Ͻg н� нH н� н)н� нM нP   P   " н3 н��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ&�Ͻ��Ͻ��Ͻ��Ͻ+ н н��Ͻ  н��Ͻ��ϽP   P   L�Ͻ��Ͻ9�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽH�Ͻ��Ͻq�Ͻ��Ͻ}�Ͻ��ϽP   P   ��Ͻ��Ͻ<�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻq�Ͻ]�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ/�Ͻ��Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ<�Ͻ9�Ͻ��Ͻ��Ͻ��Ͻ н��Ͻ
 н��Ͻ��Ͻ��ϽR�ϽR�Ͻ��Ͻ��Ͻ��Ͻa�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ3 нl нO нt н� н� н� н нE н н��Ͻ��Ͻ��Ͻ��Ͻq�ϽP   P   +�Ͻ8�Ͻ��Ͻ9 н� н,н�н�н�н�н8н�н}н�н�н,н� нD н��Ͻ.�ϽP   P   .�Ͻm�Ͻ��Ͻ& н� н н�н�нCнHн�н�н�нн�н�н�н� н н��ϽP   P   ��Ͻ �Ͻ��Ͻ8 н� н�н�н�н�нLнн�н�нAн�н�н�н�н� н нP   P   D н��Ͻ��Ͻw н� н�н�нHнQнн�нxн�н�нCн&н6н�н�н� нP   P   � н� н н н� нннн^н�н.н~н�н�н
н�нPн6н�н�нP   P   ,н� нI нn нy н;н�ннOн�нн?н�н�нYнн�н&н�н�нP   P   �нн� нp н� н� нн�н�н�н.нNн�н<	н�нYн
нCн�н�нP   P   �н� н� н� н� н� н� н�ннiн�н{н�н#	н<	н�н�н�нAннP   P   }н�н� н� н� нs н� н�н�нjн�н�н�н�н�н�н�н�н�н�нP   P   �нdн�н� нO нV н� н�нiн�н�н�н�н{нNн?н~нxн�н�нP   P   8н�н�нн^ н��Ͻf нн�н�нkн�н�н�н.нн.н�нн�нP   P   �н�н|н� н& н��Ͻ��Ͻ2 н� н�н�н�нjнiн�н�н�ннLнHнP   P   �нн�н� н��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ� н�нiн�нн�нOн^нQн�нCнP   P   �н�н�н� н/ н��Ͻ��Ͻ��Ͻ��Ͻ2 нн�н�н�н�нннHн�н�нP   P   �нн� н� н� н��Ͻ��Ͻ��Ͻ��Ͻ��Ͻf н� н� н� нн�нн�н�н�нP   P   ,нн� нk н^ н��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽV нs н� н� н;нн�н�н нP   P   � н� н� н� н� н^ н� н/ н��Ͻ& н^ нO н� н� н� нy н� н� н� н� нP   P   9 н� н_ н� н� нk н� н� н� н� нн� н� н� нp нn н нw н8 н& нP   P   ��Ͻ��Ͻ н_ н� н� н� н�н�н|н�н�н� н� н� нI н н��Ͻ��Ͻ��ϽP   P   8�Ͻ'�Ͻ��Ͻ� н� ннн�нн�н�нdн�н� нн� н� н��Ͻ �Ͻm�ϽP   P   ��Ͻ6 н� н н?н1н5н�нIн�нiн�нн�ннDн�нн� н5 нP   P   5 нk нk н-н�н�н�н�н�н�н�н�нн�нн�н�нн8н� нP   P   � н� н� нCн�нnн�н�н�н�н�нlн�н�нuн�нLнfнн8нP   P   н
н� н=н�н\н�нvн�нX	н
н�
н�
нN
н	н�н�н�нfннP   P   �н�н� н�нн�н�н�нн+	н�
н�нUн�н�
нK	н�н�нLн�нP   P   Dнн� н9н�нTнeн�н�н:	нBн�н�н�н>н�
нK	н�н�н�нP   P   н�н�н�н�н�нBн�н�нz	н�
нн�н_н�н>н�
н	нuннP   P   �н-нAн�н�н`нн�нxн�нz
н�н�нн_н�н�нN
н�н�нP   P   н�н�н,нBн?нн~нHнн�н�
нVн�н�н�нUн�
н�ннP   P   �нн�н�нdнvн�н н н�н�нXн�
н�нн�н�н�
нlн�нP   P   iнн�н�нOн� нsн�н�н н�н�н�нz
н�
нBн�
н
н�н�нP   P   �н�н�н.н<нн� нbн)н�н н�нн�нz	н:	н+	нX	н�н�нP   P   Iн$н�н:нYн� н< н� нHн)н�н нHнxн�н�нн�н�н�нP   P   �нrн�нxн]нx н��Ͻ н� нbн�н н~н�н�н�н�нvн�н�нP   P   5н н*н�н�н� н� н��Ͻ< н� нsн�нннBнeн�н�н�н�нP   P   1ннQн%нrн� н� нx н� нн� нvн?н`н�нTн�н\нnн�нP   P   ?н�н�н�н�нrн�н]нYн<нOнdнBн�н�н�нн�н�н�нP   P    н�нн�н�н%н�нxн:н.н�н�н,н�н�н9н�н=нCн-нP   P   � н� ннн�нQн*н�н�н�н�н�н�нAн�н� н� н� н� нk нP   P   6 н� н� н�н�нн нrн$н�ннн�н-н�нн�н
н� нk нP   P   � н� н� ннpн8нYн�ннgн�н�н�нOннMн�н�н� н� нP   P   � н� н� н�н@н=нPн�н 	н�
н�
н�
н�
нG	н�н.нtнkнн� нP   P   � нw н� н&нxннFн�нJ
н}н�нн�нн�	н�н�н�н>ннP   P   �н*н4н�нYн�нDн8	н�н�н�н�н|н�н�н�н^	нYн�нkнP   P   �нн�н нн�н#н�	н�н�нrн[н-н<нZн�нdн^	н�нtнP   P   Mн:н�н�н(н?н3н�нVн�нaн�нzн�нн/н�н�н�н.нP   P   н�н�нPн�н�н)н�н6
н�нAн
нJн�нннZн�н�	н�нP   P   OнWнIнnнTн=нEн�н	н<н�н>н�нRн�н�н<н�ннG	нP   P   �ннGнDн�нaнPн�н�н�
н�н�н&н�нJнzн-н|н�н�
нP   P   �н�н�н5н@нMн�н�н�нqн�
нн�н>н
н�н[н�нн�
нP   P   �н�н�н�н�нRн�н�н�н�н�н�
н�н�нAнaнrн�н�н�
нP   P   gн�н�н�нWн�н9н�н�н�н�нqн�
н<н�н�н�н�н}н�
нP   P   н|н�н�н�нн� нн�н�н�н�н�н	н6
нVн�н�нJ
н 	нP   P   �н�н�н�н�нн� нLнн�н�н�н�н�н�н�н�	н8	н�н�нP   P   Yн0н�н�н�н)нOн� н� н9н�н�нPнEн)н3н#нDнFнPнP   P   8н�нFнSн)н�н)ннн�нRнMнaн=н�н?н�н�нн=нP   P   pн9н�нVн�н)н�н�н�нWн�н@н�нTн�н(ннYнxн@нP   P   н�н�нWнVнSн�н�н�н�н�н5нDнnнPн�н н�н&н�нP   P   � н1н&н�н�нFн�н�н�н�н�н�нGнIн�н�н�н4н� н� нP   P   � н` н1н�н9н�н0н�н|н�н�н�ннWн�н:нн*нw н� нP   P   ��ϽN нBн�н6н�н�н�	н
н�
н^н�
н�	нd	н�н�н�н�нNнT нP   P   T н нkннн�н�н^
нн�н�н�н�нUнk
нmнн	нн?нP   P   Nн� нYнн�н�н%	нgн�н�н�нjнxн�н�нYн�н=н�ннP   P   �н�н�нlн?н=н�нн�нн�нн�н�н�н�нн�н=н	нP   P   �нн�нн�нн�нbн�н�н,н}н"нsнн�нlнн�ннP   P   �нhн�нmн�н�н�н^нVн�нPн нSн~н&нIн�н�нYнmнP   P   �н�нXн�н\н�н�нm
н�нWнн/н(нeнн&нн�н�нk
нP   P   d	нiнCн&н>н5н{нx	нAн�н�н�нhнUнeн~нsн�н�нUнP   P   �	нpн�нннн�нvн�	н�нuн ннhн(нSн"н�нxн�нP   P   �
н�нsн�ннн�н�н�н�
н�нQн н�н/н н}ннjн�нP   P   ^ннyнCнDнNн0н3нTнaнCн�нuн�ннPн,н�н�н�нP   P   �
н�н0н�н8нtнQн^н�ннaн�
н�н�нWн�н�нн�н�нP   P   
н�н^н�н�н� н( н� нFн�нTн�н�	нAн�нVн�н�н�ннP   P   �	н�н�нxнXн� нI н~ н� н^н3н�нvнx	нm
н^нbннgн^
нP   P   �н\н�нqнAн7нn нI н( нQн0н�н�н{н�н�н�н�н%	н�нP   P   �н�нEнHн�н�н7н� н� нtнNннн5н�н�нн=н�н�нP   P   6н�н�н,нXн�нAнXн�н8нDннн>н\н�н�н?н�ннP   P   �н�н�н�н,нHнqнxн�н�нCн�нн&н�нmннlнннP   P   Bн�нRн�н�нEн�н�н^н0нyнsн�нCнXн�н�н�нYнkнP   P   N н� н�н�н�н�н\н�н�н�нн�нpнiн�нhнн�н� н нP   P    �Ͻ]�Ͻ н�н2нyн�нG
н}н5нZн>н�нF
н�нPнHн�н* нN�ϽP   P   N�ϽG�Ͻ) нн@н�н�	н�н]нeн`нyн@н6н\н�	н�нн�н нP   P   * н��Ͻ7 н�н�н�н�
н;н�нRнZн�нLнlн�н'н�
н�н�н�нP   P   �н� н� н�нdн�н{н н�н�н�н-ннxн�н�н�нnн�ннP   P   HнMн�нWн5н�н�
н'нн�нн�н�н�нн�нн�н�
н�нP   P   Pн�н�нlннaн�	нEн�н�н#н�нн�н~н"н�н�н'н�	нP   P   �нbн�н�н�нLн�н]н�н�нн�н�н н�н~нн�н�н\нP   P   F
н�н9нн=нBн�нD
нEнbнaнн�нC н н�н�нxнlн6нP   P   �н�н{н"нн�нzн�н�нJнtн,н�н�н�нн�ннLн@нP   P   >нs	ннн�н�н]н�нp	н!нnн�н,нн�н�н�н-н�нyнP   P   Zн�	нMн+н�нpн�н%нUн
нvнnнtнaнн#нн�нZн`нP   P   5н$
н�н�н�нz н� н�н�н�н
н!нJнbн�н�н�н�нRнeнP   P   }нs	н2н�н.н� н1 н� нн�нUнp	н�нEн�н�нн�н�н]нP   P   G
н�н&нOн�н� н��Ͻ��Ͻ� н�н%н�н�нD
н]нEн'н н;н�нP   P   �н(нVнUн�н� н# н��Ͻ1 н� н�н]нzн�н�н�	н�
н{н�
н�	нP   P   yнkнcнCн�н�н� н� н� нz нpн�н�нBнLнaн�н�н�н�нP   P   2нн�нFн�н�н�н�н.н�н�н�нн=н�нн5нdн�н@нP   P   �нmн�н�нFнCнUнOн�н�н+нн"нн�нlнWн�н�ннP   P    н� н�н�н�нcнVн&н2н�нMнн{н9н�н�н�н� н7 н) нP   P   ]�Ͻ��Ͻ� нmннkн(н�нs	н$
н�	нs	н�н�нbн�нMн� н��ϽG�ϽP   P   �Ͻ#�Ͻ��Ͻ.н�ннv
н(н]н�нн�нrнUн|
н�н�нн��Ͻ#�ϽP   P   #�ϽT�ϽL�Ͻfн�ннaн�нiнBнsнOнNн�нSнLн-н�ннK�ϽP   P   ��Ͻ"�Ͻ��Ͻнн,н�н�н�н\н�н�н�нxн�н�н�ннVннP   P   н`�Ͻ_�ϽCн�нMн�нOн�н,н�н!!нA!н5н�н�н�н�нн�нP   P   �н?нD нIн�нннн�н�н�!н$нJ%нK$н�!н�н�н�н�н-нP   P   �ннxн|нLннRн�н�н�н�"н&н�'н�'н�%н�"н�н�н�нLнP   P   |
н�н
н�нн�н�
нMнн�н�!н�%н�(н�)н�(н�%н�!н�н�нSнP   P   Uн�нIнн3нrн	нJнн�нBнm$н�'н7*н�)н�'нK$н5нxн�нP   P   rнs	н�н�н�н�н�нt	н�нн�н/!н1%н�'н�(н�'нJ%нA!н�нNнP   P   �н�н�нdннн�н�н�н�нPнpн/!нm$н�%н&н$н!!н�нOнP   P   н�нZн�нlнZ�Ͻ>н�н�н�н?нPн�нBн�!н�"н�!н�н�нsнP   P   �н�н�нBнkн��Ͻ1�Ͻ;нJнgн�н�нн�н�н�н�н,н\нBнP   P   ]н�нhн�нU н��Ͻ"�Ͻ��Ͻl нJн�н�н�ннн�н�н�н�нiнP   P   (н�	н�н�н_н��Ͻ��Ͻ�Ͻ��Ͻ;н�н�нt	нJнMн�ннOн�н�нP   P   v
нUнWн�н:нf�Ͻ��Ͻ��Ͻ"�Ͻ1�Ͻ>н�н�н	н�
нRнн�н�нaнP   P   н�н�ннdн'�Ͻf�Ͻ��Ͻ��Ͻ��ϽZ�Ͻн�нrн�нннMн,ннP   P   �нgн�нiнPнdн:н_нU нkнlнн�н3ннLн�н�нн�нP   P   .н�н�ннiнн�н�н�нBн�нdн�нн�н|нIнCннfнP   P   ��Ͻq�Ͻ н�н�н�нWн�нhн�нZн�н�нIн
нxнD н_�Ͻ��ϽL�ϽP   P   #�Ͻs�Ͻq�Ͻ�нgн�нUн�	н�н�н�н�нs	н�н�нн?н`�Ͻ"�ϽT�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ�н'н�
н]нн`нkн3н=нwн�
н�н�н��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��ϽKн�н>н�н�н�н[н8н�н2н1нDнUн�нe�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ~�Ͻн)	нoн�н&н�н�"нa#н�"н�н_нfнHн�ннe�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ*нH	н�н|н(нT$н(н�)н�)н�'н$н�н0н�н�н�нP   P   �н �Ͻ	�Ͻ��Ͻ�нfн�нHн�н�%н�*н�.н0н�.н+н�%н�н0нHнUнP   P   �нн��Ͻ��Ͻ<н н?н�нPн�%н�+н�1н&4н�3нt1н�+н�%н�нfнDнP   P   �
н�н�нo н�нZн�
нbнFн$н+н�1н5нw6нk5нt1н+н$н_н1нP   P   wн�нн� н� нPн�н]нfн$ н�'н�.н4н�6нw6н�3н�.н�'н�н2нP   P   =н�
н�нwн нYн�н�
н2н�н�"н�)н0н4н5н&4н0н�)н�"н�нP   P   3нuн9нFн��Ͻ�Ͻgнн�н>нVнl#н�)н�.н�1н�1н�.н�)нa#н8нP   P   kнpн"н�н��Ͻv�Ͻ��Ͻ�нн>нlнVн�"н�'н+н�+н�*н(н�"н[нP   P   `н0н�нJн;�ϽC�Ͻd�Ͻ�ϽDн�н>н>н�н$ н$н�%н�%нT$н�н�нP   P   н�н4нrн��Ͻ�Ͻ�Ͻ��Ͻ��ϽDнн�н2нfнFнPн�н(н&н�нP   P   ]н"н5н�н'�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�нн�
н]нbн�нHн|н�н�нP   P   �
н�н�н�н��Ͻ��Ͻ��Ͻ��Ͻ�Ͻd�Ͻ��Ͻgн�н�н�
н?н�н�нoн>нP   P   'н�нoн�нO�ϽI�Ͻ��Ͻ��Ͻ�ϽC�Ͻv�Ͻ�ϽYнPнZн нfнH	н)	н�нP   P   �нGн�нн��ϽO�Ͻ��Ͻ'�Ͻ��Ͻ;�Ͻ��Ͻ��Ͻ н� н�н<н�н*ннKнP   P   ��Ͻf�Ͻ��Ͻ� нн�н�н�нrнJн�нFнwн� нo н��Ͻ��Ͻ��Ͻ~�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ�нoн�н5н4н�н"н9н�нн�н��Ͻ	�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻf�ϽGн�н�н"н�н0нpнuн�
н�н�нн �Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ/�Ͻ�Ͻ� нн�нVнн'ннн�нEнIн�н� нC�Ͻ!�Ͻ��ϽP   P   ��Ͻ��Ͻ5�Ͻ6�Ͻ�н�нн�н}н&!н�"н�"н� нCн�нн�нQн$�Ͻ��ϽP   P   !�Ͻ��Ͻ�ϽZ�Ͻ�н�нCн�н�!нM(н,н�-н,н((н�!нWн�н�н�н$�ϽP   P   C�Ͻ>�Ͻ��Ͻf�Ͻyн�н�н1н�$н-н�2нV6н96н�2н�,н�$н�н�н�нQнP   P   � н��Ͻi�Ͻ��Ͻ� н�нн5н�&н0нy7нe<н	>нY<н�7н�/н�&н�н�н�нP   P   �н
 нR�ϽU�ϽC н�нн|н�$н�/н_9н�?н�Bн�Bн�?нS9н�/н�$нWннP   P   Iн.н��Ͻ�Ͻ��Ͻ1н`н�н�!н�,н�7н�?нhDн�FнuDн�?н�7н�,н�!н�нP   P   Eн�н	н��Ͻ��ϽннAн{нZ(н�2нX<н�Bн�Fн�Fн�BнY<н�2н((нCнP   P   �н�н�н��Ͻ�Ͻ��Ͻ�нн�н&!н�+нV6н(>н�BнhDн�Bн	>н96н,н� нP   P   нн�нp�Ͻ�Ͻ	�Ͻ^�Ͻ�нAнн�"н�-нV6нX<н�?н�?нe<нV6н�-н�"нP   P   нн>н��ϽF�Ͻ��Ͻ*�Ͻ' н�н)н�н�"н�+н�2н�7н_9нy7н�2н,н�"нP   P   'н4нbнm нi�Ͻ��Ͻ��ϽZ�ϽZ н�н)нн&!нZ(н�,н�/н0н-нM(н&!нP   P   н4нeн` н��Ͻc�ϽQ�Ͻ|�Ͻ��ϽZ н�нAн�н{н�!н�$н�&н�$н�!н}нP   P   VнDн�нC н]�Ͻ��Ͻ��Ͻ��Ͻ|�ϽZ�Ͻ' н�ннAн�н|н5н1н�н�нP   P   �ннн��Ͻu�Ͻ��ϽB�Ͻ��ϽQ�Ͻ��Ͻ*�Ͻ^�Ͻ�нн`ннн�нCннP   P   нNн<н�Ͻ%�Ͻ�Ͻ��Ͻ��Ͻc�Ͻ��Ͻ��Ͻ	�Ͻ��Ͻн1н�н�н�н�н�нP   P   � н< н*�Ͻ��Ͻj�Ͻ%�Ͻu�Ͻ]�Ͻ��Ͻi�ϽF�Ͻ�Ͻ�Ͻ��Ͻ��ϽC н� нyн�н�нP   P   �Ͻ�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��ϽC н` нm н��Ͻp�Ͻ��Ͻ��Ͻ�ϽU�Ͻ��Ͻf�ϽZ�Ͻ6�ϽP   P   /�Ͻ��Ͻ��Ͻ��Ͻ*�Ͻ<нн�нeнbн>н�н�н	н��ϽR�Ͻi�Ͻ��Ͻ�Ͻ5�ϽP   P   ��Ͻ��Ͻ��Ͻ�Ͻ< нNннDн4н4ннн�н�н.н
 н��Ͻ>�Ͻ��Ͻ��ϽP   P   P�Ͻ��Ͻ��ϽJ�ϽW�Ͻ�нcнSнн�нUн�н�н�н�нsн��Ͻ��Ͻ_�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻvн%н�н�"н�(н&,н,нs(н�"н�н�н;н��Ͻ��Ͻd�ϽP   P   _�Ͻ��Ͻf�Ͻ��Ͻ��Ͻ	н�н�н�*н�2н�7н�9н|7н>2н>*нrнн�н�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�нhн"н�.н�9н�Aн�Eн�Eн�Aн�9н�.н�!нн�н��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�нPн;"н�0н�=н�Gн?Nн%Pн�Mн�Gнn=нq0н�!нн;нP   P   sн��Ͻ�Ͻ5�Ͻ��Ͻ�н"н�н/н�=н�Iн?Rн�Wн�WнLRн�Iнn=н�.нrн�нP   P   �н�н��Ͻ��Ͻ��Ͻ�н�нн`*н:н�GнrRн�Yн�\н�YнLRн�Gн�9н>*н�нP   P   �нjн��Ͻe�Ͻ>�Ͻ��Ͻ�н
н�"нa2н�Aн�Mн�Wн�\н�\н�Wн�Mн�Aн>2н�"нP   P   �н�нн	�Ͻo�Ͻ[�Ͻн�н�н�(нw7н�EнTPн�Wн�Yн�Wн%Pн�Eн|7нs(нP   P   �н�н.н�Ͻ��Ͻ~�Ͻ�Ͻ]н�н�н&,н':н�Eн�MнrRн?Rн?Nн�Eн�9н,нP   P   Uн\нн��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ�н�н1н&,нw7н�Aн�Gн�Iн�Gн�Aн�7н&,нP   P   �н�нн��Ͻ��Ͻ��Ͻr�Ͻ��Ͻ��ϽDн�н�н�(нa2н:н�=н�=н�9н�2н�(нP   P   н�ннu�Ͻ��Ͻf�Ͻ��Ͻ_�Ͻu�Ͻ��Ͻ�н�н�н�"н`*н/н�0н�.н�*н�"нP   P   Sн�н6н�Ͻ��Ͻ��Ͻy�Ͻ��Ͻ_�Ͻ��Ͻ��Ͻ]н�н
нн�н;"н"н�н�нP   P   cн�н�н9�ϽH�Ͻu�Ͻ��Ͻy�Ͻ��Ͻr�Ͻ�Ͻ�Ͻн�н�н"нPнhн�н%нP   P   �н�н��ϽI�Ͻ��ϽL�Ͻu�Ͻ��Ͻf�Ͻ��Ͻ��Ͻ~�Ͻ[�Ͻ��Ͻ�н�н�н�н	нvнP   P   W�Ͻ��Ͻ��Ͻ��Ͻ*�Ͻ��ϽH�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻo�Ͻ>�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   J�Ͻ��Ͻq�Ͻ��Ͻ��ϽI�Ͻ9�Ͻ�Ͻu�Ͻ��Ͻ��Ͻ�Ͻ	�Ͻe�Ͻ��Ͻ5�Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ�Ͻl�Ͻq�Ͻ��Ͻ��Ͻ�н6нннн.нн��Ͻ��Ͻ�Ͻ��Ͻ��Ͻf�Ͻ��ϽP   P   ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�н�н�н�н�н\н�н�нjн�н��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   |�Ͻ��Ͻ��Ͻ�ϽE�Ͻ�нFнFнDн#н %н.#н�н�н�н�нk�Ͻ��Ͻ�Ͻq�ϽP   P   q�Ͻ��Ͻ��Ͻ�ϽR�Ͻ�н�нkн+н�2нU7н7н�2н+н9нн\нJ�Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻh�Ͻ��Ͻ��Ͻ�н1нr&н�4н�@н{GнQIнXGн6@н74н&н�н�н-�Ͻ��ϽP   P   ��Ͻ*�Ͻ�Ͻ��ϽO�Ͻ�н�н;*н�;нYIнYTн�Yн�YнHTнOIнF;н�)н�н�нJ�ϽP   P   k�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ннG*н�=нsNн�\н�eн@hн_eн!\нENн�<н�)н�н\нP   P   �нe�Ͻ��Ͻ�Ͻ6�Ͻ�нmнQ&нe;нaNнp_н�kнrн(rн�kн_нENнF;н&ннP   P   �н��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�нPн�4нIнu\н�kн�uн�wн/uн�kн!\нOIн74н9нP   P   �нSн��Ͻ��ϽF�Ͻ��Ͻ\нн+н1@нtTнueн7rн�wн�wн(rн_eнHTн6@н+нP   P   �н�н=�Ͻ��Ͻ�Ͻ��ϽQ�Ͻ�н�н�2н�Gн�Yн�hн7rн�uнrн@hн�YнXGн�2нP   P   .#н�нн�Ͻ��Ͻ��Ͻ��Ͻ[нtнC#н7н^Iн�Yнueн�kн�kн�eн�YнQIн7нP   P    %нн�н��ϽG�Ͻ+�Ͻ{�Ͻ��Ͻ�нн
%н7н�GнtTнu\нp_н�\нYTн{GнU7нP   P   #н?н�н��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ннC#н�2н1@нIнaNнsNнYIн�@н�2нP   P   Dн�н�н��Ͻ�Ͻ��Ͻ �Ͻ��Ͻ�Ͻ��Ͻ�нtн�н+н�4нe;н�=н�;н�4н+нP   P   Fн�нXн��Ͻ�Ͻ��Ͻ~�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ[н�ннPнQ&нG*н;*нr&нkнP   P   Fн�н��ϽX�Ͻ�Ͻ��Ͻ4�Ͻ~�Ͻ �Ͻ��Ͻ{�Ͻ��ϽQ�Ͻ\н�нmнн�н1н�нP   P   �н$�Ͻ7�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ+�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�н�н�н�н�нP   P   E�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��ϽG�Ͻ��Ͻ�ϽF�Ͻ�Ͻ6�Ͻ��ϽO�Ͻ��ϽR�ϽP   P   �Ͻ"�ϽH�ϽL�Ͻ��Ͻ��ϽX�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   ��ϽZ�ϽM�ϽH�Ͻ��Ͻ7�Ͻ��ϽXн�н�н�нн=�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻh�Ͻ��ϽP   P   ��Ͻ��ϽZ�Ͻ"�Ͻ��Ͻ$�Ͻ�н�н�н?нн�н�нSн��Ͻe�Ͻ��Ͻ*�Ͻ��Ͻ��ϽP   P   ��Ͻ{�Ͻi�Ͻ��Ͻh�ϽO�Ͻ�ннj$н�*н-нz*н�#нKнPн��Ͻ��Ͻ�Ͻ��ϽQ�ϽP   P   Q�Ͻo�Ͻ4�Ͻ��Ͻ�Ͻ�н�н�&н*5н�?н�Eн4Eн�?н�4н4&н�нQн��ϽV�Ͻ.�ϽP   P   ��Ͻ��ϽT�Ͻ��Ͻ�Ͻkн�н�/нhBн�Qн�[н_н�[н]Qн�Aн8/н(н�нU�ϽV�ϽP   P   �ϽG�Ͻ �Ͻf�Ͻ��Ͻ^н7н�3н3Kн�^нmн%uн<uн�lнo^н�JнW3н�н�н��ϽP   P   ��Ͻ�Ͻ9�Ͻ:�Ͻ/�Ͻ�н�н�3н�Mнfн�xнÄн
�н{�н�xн�eн'MнW3н(нQнP   P   ��ϽM�Ͻ��Ͻ��Ͻ.�Ͻ"�Ͻ=н�/нKн4fн}н��нO�нP�н��н�|н�eн�Jн8/н�нP   P   Pн��Ͻ��Ͻ��Ͻ7�Ͻ_�Ͻ�н2&н�Bн�^н�xн��нQ�н[�н�н��н�xнo^н�Aн4&нP   P   Kнн��Ͻ��Ͻ��Ͻ��Ͻ�н�н5нyQнmн��н`�н�н[�нP�н{�н�lн]Qн�4нP   P   �#н�
н��Ͻ�Ͻ��ϽC�Ͻ#�Ͻ�
н2$н�?н(\н/uнU�н`�нQ�нO�н
�н<uн�[н�?нP   P   z*н;н��Ͻ�Ͻ:�Ͻ�Ͻ��Ͻ��Ͻ&н�*нUEн_н/uн��н��н��нÄн%uн_н4EнP   P   -нwн_�Ͻo�Ͻ��Ͻ�Ͻ��Ͻ=�Ͻ��ϽXн-нUEн(\нmн�xн}н�xнmн�[н�EнP   P   �*нhн4�Ͻ��Ͻ��Ͻ��Ͻm�Ͻv�Ͻ��Ͻ�ϽXн�*н�?нyQн�^н4fнfн�^н�Qн�?нP   P   j$н�н��Ͻ��Ͻ{�Ͻs�Ͻ��Ͻ;�Ͻ��Ͻ��Ͻ��Ͻ&н2$н5н�BнKн�Mн3KнhBн*5нP   P   нн�Ͻr�Ͻ��Ͻ`�Ͻ��Ͻ��Ͻ;�Ͻv�Ͻ=�Ͻ��Ͻ�
н�н2&н�/н�3н�3н�/н�&нP   P   �нsнu�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻm�Ͻ��Ͻ��Ͻ#�Ͻ�н�н=н�н7н�н�нP   P   O�Ͻ��Ͻ�Ͻv�Ͻ��Ͻd�Ͻ��Ͻ`�Ͻs�Ͻ��Ͻ�Ͻ�ϽC�Ͻ��Ͻ_�Ͻ"�Ͻ�н^нkн�нP   P   h�Ͻ��Ͻj�Ͻ.�Ͻ#�Ͻ��Ͻ��Ͻ��Ͻ{�Ͻ��Ͻ��Ͻ:�Ͻ��Ͻ��Ͻ7�Ͻ.�Ͻ/�Ͻ��Ͻ�Ͻ�ϽP   P   ��Ͻ��Ͻ/�Ͻ<�Ͻ.�Ͻv�Ͻ��Ͻr�Ͻ��Ͻ��Ͻo�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ:�Ͻf�Ͻ��Ͻ��ϽP   P   i�Ͻ|�Ͻ��Ͻ/�Ͻj�Ͻ�Ͻu�Ͻ�Ͻ��Ͻ4�Ͻ_�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ9�Ͻ �ϽT�Ͻ4�ϽP   P   {�Ͻ�Ͻ|�Ͻ��Ͻ��Ͻ��Ͻsнн�нhнwн;н�
нн��ϽM�Ͻ�ϽG�Ͻ��Ͻo�ϽP   P   G�Ͻ��Ͻl�Ͻ��ϽD�ϽG�Ͻ�
н�нV+н~4н�7н#4н+нн
н��Ͻ��Ͻ�Ͻ��Ͻ:�ϽP   P   :�Ͻ8�Ͻ�Ͻ,�Ͻ�Ͻc�Ͻ#н�-н�Aн�Pн�XнgXнgPн<Aн�,н>н��ϽS�Ͻ��Ͻ#�ϽP   P   ��Ͻ;�Ͻg�Ͻ��Ͻ��Ͻf нн�9нvTнTiнTvн�zн2vн�hнTн�8н}н��Ͻ�Ͻ��ϽP   P   �Ͻ��Ͻ��ϽF�Ͻ��Ͻb н� н�@н `н�{н4�н�н�н�н�zн\_н@н�н��ϽS�ϽP   P   ��Ͻ4�Ͻ��Ͻ��Ͻ!�Ͻ�Ͻ	н�@нkdн��нŝн$�н��н�нt�нi�н�cн@н}н��ϽP   P   ��Ͻ�Ͻ��Ͻ}�Ͻ �Ͻ��Ͻ�н|9н`н��нG�н��н:�н4�н0�н�нi�н\_н�8н>нP   P   
н�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�
нS-нzTнT{нНн~�н9�н�н	�н0�нt�н�zнTн�,нP   P   нZ�Ͻf�Ͻ�ϽB�ϽW�Ͻv�Ͻ|н�Aн3iн@�н/�нY�н(�н�н4�н�н�н�hн<AнP   P   +н�н��Ͻ��Ͻ�Ͻ�Ͻ!�Ͻ:	н,+н�Pнsvн�нϳнY�н9�н:�н��н�н2vнgPнP   P   #4н�н3�Ͻ?�ϽO�Ͻ/�ϽR�Ͻ!�Ͻ�нs4н�Xн{н�н/�н~�н��н$�н�н�zнgXнP   P   �7н�н^�Ͻ��Ͻ��Ͻ$�Ͻ!�Ͻ��Ͻ��Ͻ�нw7н�Xнsvн@�нНнG�нŝн4�нTvн�XнP   P   ~4н�н5�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�нs4н�Pн3iнT{н��н��н�{нTiн�PнP   P   V+н�н��Ͻ��Ͻ�Ͻ��Ͻ��Ͻl�Ͻ�Ͻ��Ͻ��Ͻ�н,+н�AнzTн`нkdн `нvTн�AнP   P   �н�	н��Ͻ(�ϽN�Ͻ��Ͻ�Ͻ!�Ͻl�Ͻ��Ͻ��Ͻ!�Ͻ:	н|нS-н|9н�@н�@н�9н�-нP   P   �
н�ϽK�Ͻ��Ͻz�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ!�ϽR�Ͻ!�Ͻv�Ͻ�
н�н	н� нн#нP   P   G�Ͻ�Ͻ�Ͻ��Ͻ��Ͻs�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ$�Ͻ/�Ͻ�ϽW�Ͻ��Ͻ��Ͻ�Ͻb нf нc�ϽP   P   D�Ͻ��Ͻ4�Ͻ��Ͻ�Ͻ��Ͻz�ϽN�Ͻ�Ͻ�Ͻ��ϽO�Ͻ�ϽB�Ͻ��Ͻ �Ͻ!�Ͻ��Ͻ��Ͻ�ϽP   P   ��Ͻ�Ͻ.�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ(�Ͻ��Ͻ��Ͻ��Ͻ?�Ͻ��Ͻ�Ͻ��Ͻ}�Ͻ��ϽF�Ͻ��Ͻ,�ϽP   P   l�ϽJ�Ͻ��Ͻ.�Ͻ4�Ͻ�ϽK�Ͻ��Ͻ��Ͻ5�Ͻ^�Ͻ3�Ͻ��Ͻf�Ͻ��Ͻ��Ͻ��Ͻ��Ͻg�Ͻ�ϽP   P   ��Ͻ��ϽJ�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ�	н�н�н�н�н�нZ�Ͻ�Ͻ�Ͻ4�Ͻ��Ͻ;�Ͻ8�ϽP   P   ȘϽm�Ͻ��Ͻ`�ϽY�Ͻ��Ͻ6	н!н�3н�?н�Cн=?нK3нE н�нz�Ͻ��Ͻ��Ͻ�Ͻ�ϽP   P   �Ͻ��ϽŦϽT�Ͻ��ϽD�Ͻ�нi8нgSнFgнqн=qн�fн�Rн=7н�н�Ͻ��Ͻ��Ͻ4�ϽP   P   �Ͻ��Ͻe�ϽL�Ͻm�Ͻ\�Ͻ� н{Hн�kн��н�н��н,�нG�н�kнmGн= нd�Ͻ��Ͻ��ϽP   P   ��ϽR�Ͻ��ϽźϽ{�ϽI�Ͻ�#н�Pн�{н�н��н�н��н��н�н�zн�Oн�"нd�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ7�Ͻ
�Ͻ��Ͻ� н�Pнz�н�нq�н��нw�н��н��н��н�н�Oн= н�ϽP   P   z�Ͻ%�Ͻ��Ͻt�Ͻ��Ͻ��Ͻ�нOHн�{н�н�н��нKѽMѽ�н��н��н�zнmGн�нP   P   �н��Ͻ��Ͻ��Ͻ��ϽO�Ͻ�н8н�kн��н��н��нnѽ�ѽ~ѽ�н��н�н�kн=7нP   P   E н]�Ͻ �Ͻ)�Ͻ��Ͻ�Ͻ��Ͻ� н<Sн&�н�н��нmѽ�ѽ�ѽMѽ��н��нG�н�RнP   P   K3нtнO�Ͻ]�Ͻ��Ͻe�Ͻ|�ϽнN3н
gнC�н�н��нmѽnѽKѽw�н��н,�н�fнP   P   =?н
н'�Ͻb�Ͻz�Ͻj�Ͻ��Ͻ �ϽTн�?н_qнԠн�н��н��н��н��н�н��н=qнP   P   �Cн�н#�Ͻ��Ͻ�Ͻq�Ͻ�Ͻ��Ͻ;�Ͻ�н�Cн_qнC�н�н��н�нq�н��н�нqнP   P   �?н�нi�Ͻ}�Ͻ��Ͻ6�ϽK�Ͻ��Ͻy�Ͻ:�Ͻ�н�?н
gн&�н��н�н�н�н��нFgнP   P   �3нWн�Ͻ��ϽJ�ϽާϽ�Ͻ֧Ͻ�Ͻy�Ͻ;�ϽTнN3н<Sн�kн�{нz�н�{н�kнgSнP   P   !н�н��Ͻ�ϽиϽ�Ͻ�ϽȟϽ֧Ͻ��Ͻ��Ͻ �Ͻн� н8нOHн�Pн�Pн{Hнi8нP   P   6	нa�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�ϽK�Ͻ�Ͻ��Ͻ|�Ͻ��Ͻ�н�н� н�#н� н�нP   P   ��Ͻ��Ͻ��Ͻ��Ͻ�ϽϳϽ��Ͻ�ϽާϽ6�Ͻq�Ͻj�Ͻe�Ͻ�ϽO�Ͻ��Ͻ��ϽI�Ͻ\�ϽD�ϽP   P   Y�ϽT�Ͻ��Ͻ(�Ͻ:�Ͻ�Ͻ��ϽиϽJ�Ͻ��Ͻ�Ͻz�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ
�Ͻ{�Ͻm�Ͻ��ϽP   P   `�ϽԽϽe�Ͻ��Ͻ(�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ}�Ͻ��Ͻb�Ͻ]�Ͻ)�Ͻ��Ͻt�Ͻ7�ϽźϽL�ϽT�ϽP   P   ��Ͻ0�Ͻ3�Ͻe�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻi�Ͻ#�Ͻ'�ϽO�Ͻ �Ͻ��Ͻ��Ͻ��Ͻ��Ͻe�ϽŦϽP   P   m�ϽĢϽ0�ϽԽϽT�Ͻ��Ͻa�Ͻ�нWн�н�н
нtн]�Ͻ��Ͻ%�Ͻ��ϽR�Ͻ��Ͻ��ϽP   P   glϽcrϽ�Ͻg�Ͻe�ϽU�ϽYн%н)?нxPн$Vн�Oн�>н$н(н��Ͻw�Ͻl�Ͻ��Ͻ�qϽP   P   �qϽ!rϽ�Ͻ��Ͻ��Ͻ��Ͻ�н�Cнiiн��н[�н��н�н7hнHBнfнh�Ͻ�Ͻ��Ͻ�~ϽP   P   ��ϽCzϽ\�Ͻ��Ͻ��Ͻ��Ͻ�%н5[н��н�н��н��н��н0�н؉н�Yн�$н��Ͻ�Ͻ��ϽP   P   l�ϽʈϽ	�Ͻ�Ͻ�Ͻ��Ͻ0*н�fн̠н7�нH�н�ѽnѽ��н9�н��н�eн�(н��Ͻ�ϽP   P   w�Ͻ�ϽʓϽb�Ͻ�Ͻ��Ͻ�%н�fн��н��нhѽL0ѽ�:ѽ0ѽ�ѽ��н̦н�eн�$нh�ϽP   P   ��Ͻ5�Ͻi�ϽZ�Ͻ޶Ͻ��Ͻwн[н�н��н�ѽ'EѽU[ѽ[ѽhDѽ,ѽ��н��н�YнfнP   P   (н�Ͻ5�ϽϥϽ[�Ͻ��Ͻ�нiCнL�н��нiѽEѽafѽtrѽNfѽhDѽ�ѽ9�н؉нHBнP   P   $н��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ@�Ͻ�$нiнE�нW�н�0ѽt[ѽ�rѽtrѽ[ѽ0ѽ��н0�н7hнP   P   �>нA�Ͻ��ϽM�Ͻ!�ϽX�Ͻ��Ͻ��Ͻ�>н��нU�н	ѽ;ѽt[ѽafѽU[ѽ�:ѽnѽ��н�нP   P   �Oн�нt�ϽB�Ͻ�Ͻ �ϽĳϽ~�Ͻ#н$PнǒнN�н	ѽ�0ѽEѽ'EѽL0ѽ�ѽ��н��нP   P   $Vн@н��Ͻ"�Ͻ�Ͻv�Ͻ��ϽG�Ͻ��ϽDн5VнǒнU�нW�нiѽ�ѽhѽH�н��н[�нP   P   xPн]нh�Ͻ�Ͻ_�Ͻi�Ͻ��ϽQ�ϽطϽN�ϽDн$Pн��нE�н��н��н��н7�н�н��нP   P   )?н-н�Ͻ!�Ͻ��Ͻ"�Ͻv{Ͻ�Ͻ`�ϽطϽ��Ͻ#н�>нiнL�н�н��н̠н��нiiнP   P   %н� нB�Ͻ��Ͻ��Ͻd�Ͻ�vϽUvϽ�ϽQ�ϽG�Ͻ~�Ͻ��Ͻ�$нiCн[н�fн�fн5[н�CнP   P   Yн��Ͻs�Ͻ&�Ͻ��Ͻ�Ͻ~{Ͻ�vϽv{Ͻ��Ͻ��ϽųϽ��Ͻ@�Ͻ�нwн�%н0*н�%н�нP   P   U�Ͻa�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ�Ͻd�Ͻ"�Ͻi�Ͻv�Ͻ �ϽX�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   e�Ͻ��Ͻp�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ_�Ͻ�Ͻ�Ͻ!�Ͻ�Ͻ[�Ͻ޶Ͻ�Ͻ�Ͻ��Ͻ��ϽP   P   g�ϽV�Ͻx�Ͻ�Ͻ��Ͻ��Ͻ&�Ͻ��Ͻ!�Ͻ�Ͻ"�ϽB�ϽM�Ͻ��ϽϥϽZ�Ͻb�Ͻ�Ͻ��Ͻ��ϽP   P   �ϽΉϽ��Ͻx�Ͻp�Ͻ�Ͻs�ϽB�Ͻ�Ͻh�Ͻ��Ͻt�Ͻ��Ͻ��Ͻ5�Ͻi�ϽʓϽ	�Ͻ\�Ͻ�ϽP   P   crϽ�zϽΉϽV�Ͻ��Ͻa�Ͻ��Ͻ� н-н]н@н�нA�Ͻ��Ͻ�Ͻ5�Ͻ�ϽʈϽCzϽ!rϽP   P   �/Ͻo8Ͻ�NϽkqϽ:�Ͻ��Ͻ��Ͻ�*н�Mн�cнSjн�bн�Lнq)н��Ͻ��Ͻ��Ͻ�oϽ�MϽ�7ϽP   P   �7Ͻ�8Ͻ�KϽ�nϽ�Ͻ��Ͻ�н�Tнۆн!�н��нZ�н|�нd�нSн�н��Ͻ!�Ͻ�mϽ6KϽP   P   �MϽ�AϽ)NϽ�nϽ�ϽW�Ͻn*н�rн��н��н�	ѽѽB	ѽ��н�нCqн�(н��Ͻh�Ͻ�mϽP   P   �oϽ�VϽ�VϽqϽ9�ϽC�Ͻf0нB�н��н^ѽFѽT_ѽ9_ѽ?EѽEѽ�н��н�.н��Ͻ!�ϽP   P   ��ϽsϽPeϽusϽY�Ͻ(�Ͻ**н��н��н>,ѽjlѽ3�ѽ�ѽڕѽFkѽ�*ѽ&�н��н�(н��ϽP   P   ��Ͻ]�ϽxϽvxϽ*�Ͻ%�Ͻ�н�rн��нB,ѽ�yѽ�ѽb�ѽ��ѽ�ѽ�xѽ�*ѽ�нCqн�нP   P   ��Ͻ.�Ͻ~�Ͻa}ϽʌϽ��Ͻ��ϽKTнh�нMѽlѽ0�ѽ��ѽ��ѽ9�ѽ�ѽFkѽEѽ�нSнP   P   q)н��Ͻ��Ͻg�Ͻ��ϽI�Ͻ��Ͻ[*нD�н�н Fѽ|�ѽ��ѽ��ѽ��ѽ��ѽڕѽ?Eѽ��нd�нP   P   �Lн��Ͻ#�Ͻo�Ͻ�{Ͻ{�Ͻ��Ͻ��ϽoMн(�н
ѽ�_ѽj�ѽ��ѽ��ѽb�ѽ�ѽ9_ѽB	ѽ|�нP   P   �bнPнO�ϽӏϽrtϽ�tϽ�Ͻ��Ͻ�н^cн��н�ѽ�_ѽ|�ѽ0�ѽ�ѽ3�ѽT_ѽѽZ�нP   P   Sjн�н��ϽҔϽLoϽ�aϽHoϽєϽ�Ͻ�н�jн��н
ѽ Fѽlѽ�yѽjlѽFѽ�	ѽ��нP   P   �cн�н�Ͻ�ϽakϽ�SϽ�SϽTkϽ�Ͻ�Ͻ�н^cн(�н�нMѽB,ѽ>,ѽ^ѽ��н!�нP   P   �Mн+нs�ϽQ�Ͻ%jϽNϽ6DϽ�MϽ�iϽ�Ͻ�Ͻ�нoMнD�нh�н��н��н��н��нۆнP   P   �*н��Ͻg�Ͻ`�Ͻ�kϽ/NϽq>Ͻ9>Ͻ�MϽTkϽєϽ��Ͻ��Ͻ[*нKTн�rн��нB�н�rн�TнP   P   ��Ͻs�Ͻc�Ͻ��ϽpϽ�TϽ[DϽq>Ͻ6DϽ�SϽHoϽ�Ͻ��Ͻ��Ͻ��Ͻ�н**нf0нn*н�нP   P   ��Ͻ��ϽD�Ͻ��Ͻ�uϽ6bϽ�TϽ/NϽNϽ�SϽ�aϽ�tϽ{�ϽI�Ͻ��Ͻ%�Ͻ(�ϽC�ϽW�Ͻ��ϽP   P   :�Ͻ2�Ͻ(�Ͻ��Ͻ}Ͻ�uϽpϽ�kϽ%jϽakϽLoϽrtϽ�{Ͻ��ϽʌϽ*�ϽY�Ͻ9�Ͻ�Ͻ�ϽP   P   kqϽ�tϽ�yϽ�~Ͻ��Ͻ��Ͻ��Ͻ`�ϽQ�Ͻ�ϽҔϽӏϽo�Ͻg�Ͻa}ϽvxϽusϽqϽ�nϽ�nϽP   P   �NϽ�WϽ�fϽ�yϽ(�ϽD�Ͻc�Ͻg�Ͻs�Ͻ�Ͻ��ϽO�Ͻ#�Ͻ��Ͻ~�ϽxϽPeϽ�VϽ)NϽ�KϽP   P   o8Ͻ�BϽ�WϽ�tϽ2�Ͻ��Ͻs�Ͻ��Ͻ+н�н�нPн��Ͻ��Ͻ.�Ͻ]�ϽsϽ�VϽ�AϽ�8ϽP   P   %�ν^�ν3Ͻs5ϽWpϽ��Ͻ��Ͻ�/н�_н^н�н�~н^нv-нR�Ͻ��Ͻ�mϽ|3Ͻ�Ͻ��νP   P   ��νZ�νZϽ�3Ͻ�vϽq�Ͻ�н�iн��н��н��нG�н��н��н�gн5н3�Ͻ�tϽ�1ϽsϽP   P   �Ͻm�ν2Ͻb3ϽyϽ��Ͻ\1нΒн��н�2ѽ`ѽfoѽ:_ѽ,1ѽ~�н��н�.н��Ͻ�vϽ�1ϽP   P   |3ϽeϽ�Ͻ�4Ͻ�uϽ��Ͻ�9н��н�ѽ�nѽK�ѽ]�ѽD�ѽ�ѽ2mѽ�ѽԦнq7н��Ͻ�tϽP   P   �mϽ8Ͻ=&Ͻ�8ϽoϽ�Ͻ 1н��нU"ѽ��ѽH�ѽeҽ21ҽ�ҽ��ѽ�ѽ�ѽԦн�.н3�ϽP   P   ��Ͻ�eϽ�>ϽC?Ͻ�fϽ$�Ͻ�н��нlѽ��ѽ��ѽ�DҽOmҽ�lҽMDҽ��ѽ�ѽ�ѽ��н5нP   P   R�Ͻ��Ͻ$[Ͻ9GϽ�[Ͻo�Ͻ�Ͻiн��н�nѽV�ѽ3Eҽ��ҽ{�ҽ�ҽMDҽ��ѽ2mѽ~�н�gнP   P   v-н��ϽwϽ�OϽ�OϽxϽ��Ͻ�.н�нo2ѽ_�ѽ�ҽ�mҽo�ҽ{�ҽ�lҽ�ҽ�ѽ,1ѽ��нP   P   ^н+�Ͻ��ϽXϽ�DϽlXϽt�Ͻ��Ͻt_н��н\`ѽ�ѽ�1ҽ�mҽ��ҽOmҽ21ҽD�ѽ:_ѽ��нP   P   �~н�	н�Ͻ�_Ͻ�9Ͻ+:Ͻ�_Ͻ��Ͻc
н8н�нpѽ�ѽ�ҽ3Eҽ�Dҽeҽ]�ѽfoѽG�нP   P   �н�нδϽ�eϽ	3ϽQ"ϽI3Ͻ�eϽ�Ͻ�нu�н�н\`ѽ_�ѽV�ѽ��ѽH�ѽK�ѽ`ѽ��нP   P   ^н�н��Ͻ�hϽ:.Ͻ�Ͻ{ϽY.Ͻ�hϽ��Ͻ�н8н��нo2ѽ�nѽ��ѽ��ѽ�nѽ�2ѽ��нP   P   �_н�
н}�Ͻ:iϽY-ϽϽ��ν�Ͻ-Ͻ�hϽ�Ͻc
нt_н�н��нlѽU"ѽ�ѽ��н��нP   P   �/н}�Ͻ;�ϽgfϽ�.ϽϽ��ν��ν�ϽY.Ͻ�eϽ��Ͻ��Ͻ�.нiн��н��н��нΒн�iнP   P   ��Ͻ��ϽϽ�`Ͻ*4ϽCϽ#�ν��ν��ν{ϽI3Ͻ�_Ͻt�Ͻ��Ͻ�Ͻ�н 1н�9н\1н�нP   P   ��Ͻ�ϽSyϽ�YϽb;ϽI#ϽCϽϽϽ�ϽQ"Ͻ+:ϽlXϽxϽo�Ͻ$�Ͻ�Ͻ��Ͻ��Ͻq�ϽP   P   WpϽhϽ]]Ͻ�QϽ�FϽb;Ͻ*4Ͻ�.ϽY-Ͻ:.Ͻ	3Ͻ�9Ͻ�DϽ�OϽ�[Ͻ�fϽoϽ�uϽyϽ�vϽP   P   s5Ͻ�9Ͻ�@Ͻ IϽ�QϽ�YϽ�`ϽgfϽ:iϽ�hϽ�eϽ�_ϽXϽ�OϽ9GϽC?Ͻ�8Ͻ�4Ͻb3Ͻ�3ϽP   P   3Ͻ�Ͻ2(Ͻ�@Ͻ]]ϽSyϽϽ;�Ͻ}�Ͻ��ϽδϽ�Ͻ��ϽwϽ$[Ͻ�>Ͻ=&Ͻ�Ͻ2ϽZϽP   P   ^�ν��ν�Ͻ�9ϽhϽ�Ͻ��Ͻ}�Ͻ�
н�н�н�	н+�Ͻ��Ͻ��Ͻ�eϽ8ϽeϽm�νZ�νP   P   Xpν�~νy�ν��νM5Ͻ��Ͻ��Ͻ38н�xн�н̯н�нxvнg5нd�Ͻ܉Ͻ�1Ͻ��ν��ν�}νP   P   �}ν6~ν}�ν��ν&<Ͻ�Ͻ4н҄н�н|%ѽhHѽ�Gѽ�#ѽ�н�нн�Ͻ�9Ͻ��ν�νP   P   ��ν�ν��ν��ν�=ϽδϽ�8нj�н6ѽ�ѽ,�ѽL�ѽY�ѽI�ѽ3ѽX�нI5н��Ͻ0;Ͻ��νP   P   ��νߴν��νZ�ν�;ϽA�ϽjCн��н�lѽ��ѽ�Cҽ�rҽ�rҽ�Aҽv�ѽjѽ��н�@н��Ͻ�9ϽP   P   �1Ͻ�νY�ν��ν�3Ͻ��ϽK8н�нV~ѽmҽ�ҽ��ҽ �ҽ��ҽ�ҽ ҽ{ѽ��нI5н�ϽP   P   ܉Ͻ�%Ͻ��ν �ν'Ͻ��Ͻ5н�нPlѽ|ҽ��ҽ�ӽ:Dӽ�Cӽ�ӽ��ҽ ҽjѽX�ннP   P   d�Ͻ�fϽ'Ͻ)�νϽ/hϽ��Ͻ?�н�5ѽ��ѽ��ҽ�ӽ|`ӽ�|ӽ�_ӽ�ӽ�ҽu�ѽ3ѽ�нP   P   g5н��Ͻ=Ͻ�Ͻ�Ͻ >Ͻ	�Ͻ*7н��нߕѽ�Cҽ*�ҽ�Dӽ}ӽ�|ӽ�Cӽ��ҽ�AҽI�ѽ�нP   P   xvн��Ͻ�`Ͻ�ϽU�ν4Ͻ�aϽ�Ͻ1xн�%ѽ��ѽ�sҽ��ҽ�Dӽ|`ӽ:Dӽ �ҽ�rҽY�ѽ�#ѽP   P   �ннs}Ͻ!Ͻ/�ν��νDϽn~Ͻfн�н�Hѽ%�ѽ�sҽ*�ҽ�ӽ�ӽ��ҽ�rҽL�ѽ�GѽP   P   ̯н�н��Ͻ�%Ͻ��ν��ν�ν�%ϽސϽiн]�н�Hѽ��ѽ�Cҽ��ҽ��ҽ�ҽ�Cҽ,�ѽhHѽP   P   �нrнo�Ͻ^*Ͻ�ν�ν��νl�ν^*Ͻ_�Ͻiн�н�%ѽߕѽ��ѽ|ҽmҽ��ѽ�ѽ|%ѽP   P   �xн�н�Ͻ�*Ͻ-�νx�ν_�νL�ν��ν^*ϽސϽfн1xн��н�5ѽPlѽV~ѽ�lѽ6ѽ�нP   P   38н��Ͻ+Ͻ�&Ͻ�ν��ν.�ν[�νL�νl�ν�%Ͻn~Ͻ�Ͻ*7н?�н�н�н��нj�н҄нP   P   ��Ͻ$�ϽCcϽ�ϽU�ν`�ν+�ν.�ν_�ν��ν�νDϽ�aϽ	�Ͻ��Ͻ5нK8нjCн�8н4нP   P   ��Ͻ�iϽ�?Ͻ�Ͻ��ν1�ν`�ν��νx�ν�ν��ν��ν4Ͻ >Ͻ/hϽ��Ͻ��ϽA�ϽδϽ�ϽP   P   M5Ͻ�(Ͻ.Ͻ�Ͻ��ν��νU�ν�ν-�ν�ν��ν/�νV�ν�ϽϽ'Ͻ�3Ͻ�;Ͻ�=Ͻ&<ϽP   P   ��νQ�νK�ν��ν�Ͻ�Ͻ�Ͻ�&Ͻ�*Ͻ^*Ͻ�%Ͻ!Ͻ�Ͻ�Ͻ)�ν �ν��νZ�ν��ν��νP   P   y�ν�ν��νK�ν.Ͻ�?ϽCcϽ+Ͻ�Ͻo�Ͻ��Ͻs}Ͻ�`Ͻ=Ͻ'Ͻ��νY�ν��ν��ν}�νP   P   �~νD�ν�νQ�ν�(Ͻ�iϽ$�Ͻ��Ͻ�нrн�нн��Ͻ��Ͻ�fϽ�%Ͻ�νߴν�ν6~νP   P   ��ͽR�ͽr#ν[wν��νYϽ��Ͻ�?н�н��н��н
�нo�н<н��Ͻ�TϽ_�ν�sνB!ν�ͽP   P   �ͽm�ͽ�ν*sν��ν�|Ͻ<нa�нA&ѽ��ѽ�ѽC�ѽH�ѽt#ѽ��н�н�xϽ��ν.pνHνP   P   B!νν�"ν�rνR�ν+�Ͻ�Aн��нS�ѽ�ҽ�pҽ��ҽ{oҽrҽ��ѽz�нT=нƋϽ��ν.pνP   P   �sν�6νr7ν~uν��ν{�Ͻ~PнZѽ��ѽ��ҽ�ӽ�Hӽ!Hӽ�ӽV�ҽQ�ѽ9ѽ�LнƋϽ��νP   P   _�ν�{ν�Zν�|ν��ν�{Ͻ"Aн�ѽ��ѽ��ҽ/jӽ$�ӽC�ӽ��ӽ�gӽ��ҽ��ѽ9ѽT=н�xϽP   P   �TϽ��ν�νn�νH�ν_WϽPн�н��ѽ�ҽ��ӽ�ԽQgԽ�fԽԽ��ӽ��ҽQ�ѽz�н�нP   P   ��ϽO$Ͻ��νf�ν�ν3&Ͻr�Ͻ��н	�ѽ�ҽ2jӽԽ��Խ��Խ؍ԽԽ�gӽV�ҽ��ѽ��нP   P   <нSyϽ|�νӤν,�ν��νI{Ͻ^>н&ѽ�ҽgӽ��ӽ
hԽa�Խ��Խ�fԽ��ӽ�ӽrҽt#ѽP   P   o�н�ϽϽ&�ν�ν�ν@Ͻ��Ͻd�н��ѽ�qҽ�IӽW�ӽ
hԽ��ԽQgԽC�ӽ!Hӽ{oҽH�ѽP   P   
�н{�Ͻ�DϽ��νVν�νV�ν�EϽ��Ͻ)�н˴ѽЎҽ�Iӽ��ӽԽ�Խ$�ӽ�Hӽ��ҽC�ѽP   P   ��н�н�^Ͻ�νrνQRν4rν��ν=_Ͻ�нc�н˴ѽ�qҽgӽ2jӽ��ӽ/jӽ�ӽ�pҽ�ѽP   P   ��н�н[hϽ>�νkνy3ν`3νEkνb�νZhϽ�н)�н��ѽ�ҽ�ҽ�ҽ��ҽ��ҽ�ҽ��ѽP   P   �н6�Ͻ�_Ͻ{�ν�gν�"ν�
ν�"ν/gνb�ν=_Ͻ��Ͻd�н&ѽ	�ѽ��ѽ��ѽ��ѽS�ѽA&ѽP   P   �?н��Ͻ�FϽ��ν�kν'#ν
�ͽ�ͽ�"νEkν��ν�EϽ��Ͻ^>н��н�н�ѽZѽ��нa�нP   P   ��Ͻ�|Ͻ: Ͻ��ν�sνR4ν�ν
�ͽ�
ν`3ν4rνV�ν@ϽI{Ͻr�ϽPн"Aн~Pн�Aн<нP   P   YϽ=(Ͻ�ν �ν��νKTνR4ν'#ν�"νy3νQRν�ν�ν��ν3&Ͻ_WϽ�{Ͻ{�Ͻ+�Ͻ�|ϽP   P   ��νo�νӼν�ν�ν��ν�sν�kν�gνkνrνVν�ν,�ν�νH�ν��ν��νR�ν��νP   P   [wν�~νj�ν��ν�ν �ν��ν��ν{�ν>�ν�ν��ν&�νӤνf�νn�ν�|ν~uν�rν*sνP   P   r#ν{9ν�]νj�νӼν�ν: Ͻ�FϽ�_Ͻ[hϽ�^Ͻ�DϽϽ|�ν��ν�ν�Zνr7ν�"ν�νP   P   R�ͽ�ν{9ν�~νo�ν=(Ͻ�|Ͻ��Ͻ6�Ͻ�н�н{�Ͻ�ϽSyϽO$Ͻ��ν�{ν�6ννm�ͽP   P   �ͽ�)ͽBqͽ��ͽQqνJϽմϽMIн��н,ѽ�'ѽ�ѽl�н�Dн��Ͻ�ϽFlν��ͽLnͽ(ͽP   P   (ͽ�(ͽ{fͽ��ͽ �νBϽн��н��ѽ� ҽ�Aҽ�@ҽ��ѽ�ѽG�н\нd<Ͻ{ν�ͽ�cͽP   P   LnͽpJͽ pͽ��ͽk�ν�[Ͻ�Lнx@ѽ�ҽ.�ҽ=Dӽ'kӽrBӽ��ҽҽ�:ѽ�FнJVϽ�ν�ͽP   P   ��ͽT�ͽJ�ͽ��ͽYνO[Ͻ,aн�wѽa�ҽ�jӽxԽ~mԽ�lԽ�Խ�fӽH~ҽ�qѽ�[нJVϽ{νP   P   Flν�ͽ0�ͽ��ͽOoν�@Ͻ�Kн�wѽ�ҽ��ӽ��Խ�*ս�[ս�(ս��Խ�ӽ��ҽ�qѽ�Fнd<ϽP   P   �Ͻ�Uν{�ͽ(�ͽ2Xν1Ͻн�?ѽ�ҽɼӽ%�Խߍս��ս��սZ�ս��Խ�ӽH~ҽ�:ѽ\нP   P   ��ϽW�ν:νnνW;ν��ν�Ͻh�н�ҽ(kӽ�Խ�ս�+ֽ�bֽ�*ֽZ�ս��Խ�fӽҽG�нP   P   �Dн�=ϽU�ν�ν�ν��ν<@Ͻ=Hнm�ѽg�ҽԽ�+ս}�սdcֽ�bֽ��ս�(ս�Խ��ҽ�ѽP   P   l�нʠϽ��ν3ν�ν�3νi�ν>�Ͻ&�н� ҽ|EӽoԽR]ս}�ս�+ֽ��ս�[ս�lԽrBӽ��ѽP   P   �ѽ��Ͻ��ν.Gν��ͽ<�ͽIHν�ν��Ͻ�ѽCҽ�lӽoԽ�+ս�սߍս�*ս~mԽ'kӽ�@ҽP   P   �'ѽ>нϽ-Wν9�ͽ�ͽ}�ͽ�Wν�Ͻ�н�(ѽCҽ|EӽԽ�Խ%�Խ��ԽxԽ=Dӽ�AҽP   P   ,ѽYн\&Ͻ&`ν_�ͽ��ͽцͽu�ͽr`ν�&Ͻ�н�ѽ� ҽg�ҽ(kӽɼӽ��ӽ�jӽ.�ҽ� ҽP   P   ��нi�ϽdϽ�`ν�ͽ*qͽ+Qͽqͽ��ͽr`ν�Ͻ��Ͻ&�нm�ѽ�ҽ�ҽ�ҽa�ҽ�ҽ��ѽP   P   MIн��Ͻ}�ν_Yν��ͽ�qͽ�>ͽe>ͽqͽu�ͽ�Wν�ν>�Ͻ=Hнh�н�?ѽ�wѽ�wѽx@ѽ��нP   P   մϽTBϽy�νSJν	�ͽ�ͽ�Qͽ�>ͽ+Qͽцͽ}�ͽIHνi�ν<@Ͻ�Ͻн�Kн,aн�LннP   P   JϽZ�νӄν�6ν��ͽN�ͽ�ͽ�qͽ*qͽ��ͽ�ͽ<�ͽ�3ν��ν��ν1Ͻ�@ϽO[Ͻ�[ϽBϽP   P   Qqν[ν�>ν(!ν�ν��ͽ	�ͽ��ͽ�ͽ_�ͽ9�ͽ��ͽ�ν�νW;ν2XνOoνYνk�ν �νP   P   ��ͽ��ͽ��ͽ�ν(!ν�6νSJν_Yν�`ν&`ν-Wν.Gν3ν�νnν(�ͽ��ͽ��ͽ��ͽ��ͽP   P   Bqͽ��ͽ�ͽ��ͽ�>νӄνy�ν}�νdϽ\&ϽϽ��ν��νU�ν:ν{�ͽ0�ͽJ�ͽ pͽ{fͽP   P   �)ͽ�Lͽ��ͽ��ͽ[νZ�νTBϽ��Ͻi�ϽYн>н��ϽʠϽ�=ϽW�ν�Uν�ͽT�ͽpJͽ�(ͽP   P   ��˽�!̽��̽ͽ��ͽV�ν��Ͻ�Uн[�н�`ѽ��ѽV^ѽ9�нHPнڄϽ�ν_�ͽDͽ�}̽a̽P   P   a̽� ̽nt̽�ͽ��ͽ�ν�н�ѽ��ѽ�ҽӽ�ӽ|�ҽ��ѽ�ѽнp�ν��ͽHͽ/q̽P   P   �}̽�L̽�̽�ͽ��ͽFϽ�ZнեѽQ�ҽ��ӽ"fԽ��Խ�cԽG�ӽ8�ҽa�ѽ?Sн Ͻ�ͽHͽP   P   Dͽ(�̽&�̽�ͽ]�ͽ�Ͻcvн3�ѽ_ӽ��Խ8�ս&�ս��սb~ս�ԽXӽz�ѽ�nн Ͻ��ͽP   P   _�ͽͽ��̽L ͽJ�ͽ��ν$Zн��ѽ��ӽ
ս�:ֽ� ׽�C׽]�ֽ�6ֽ�ս��ӽz�ѽ?Sнp�νP   P   �ν�ͽe1ͽ2ͽ9�ͽԬν3н�ѽ_ӽ,
ս�zֽX�׽ؽ�ؽ�׽vֽ�սXӽa�ѽнP   P   ڄϽ{OνF�ͽ�Iͽ�ͽ�Rν��ϽPѽR�ҽ�Խ�;ֽ��׽dؽy�ؽ|bؽ�׽�6ֽ�Խ8�ҽ�ѽP   P   HPн��ν��ͽ�eͽ�fͽS�ͽ'�ν�Tн3�ѽ��ӽ�ս ׽*ؽ��ؽy�ؽ�ؽ]�ֽb~սG�ӽ��ѽP   P   8�н�pϽ�Bν��ͽCͽ��ͽEEνtϽ�н`�ҽ�gԽf�սCF׽*ؽdؽؽ�C׽��ս�cԽ|�ҽP   P   V^ѽm�Ͻ��ν��ͽ}$ͽ�$ͽ�ͽ��ν�Ͻ�aѽ�ӽJ�Խf�ս ׽��׽X�׽� ׽&�ս��Խ�ӽP   P   ��ѽ�
н4�ν��ͽqͽ	�̽�ͽȶͽ�ν нx�ѽ�ӽ�gԽ�ս�;ֽ�zֽ�:ֽ8�ս"fԽӽP   P   �`ѽlн��νC�ͽFͽK�̽��̽/ͽ��ͽY�ν н�aѽ`�ҽ��ӽ�Խ,
ս
ս��Խ��ӽ�ҽP   P   [�н��Ͻ�νM�ͽ�̽��̽�W̽s�̽&�̽��ͽ�ν�Ͻ�н3�ѽR�ҽ_ӽ��ӽ_ӽQ�ҽ��ѽP   P   �Uн�uϽE�ν�ͽ�ͽ*�̽7@̽�?̽s�̽/ͽȶͽ��νtϽ�TнPѽ�ѽ��ѽ3�ѽեѽ�ѽP   P   ��Ͻ��ν|Gν��ͽ�ͽ[�̽:X̽7@̽�W̽��̽�ͽ�ͽEEν'�ν��Ͻ3н$Zнcvн�Zн�нP   P   V�νVν��ͽ��ͽc(ͽk�̽[�̽*�̽��̽K�̽	�̽�$ͽ��ͽS�ͽ�RνԬν��ν�ϽFϽ�νP   P   ��ͽ�ͽ�ͽ,kͽ�Fͽc(ͽ�ͽ�ͽ�̽Fͽqͽ}$ͽCͽ�fͽ�ͽ9�ͽJ�ͽ]�ͽ��ͽ��ͽP   P   ͽQ$ͽ27ͽ
Oͽ,kͽ��ͽ��ͽ�ͽM�ͽC�ͽ��ͽ��ͽ��ͽ�eͽ�Iͽ2ͽL ͽ�ͽ�ͽ�ͽP   P   ��̽��̽n�̽27ͽ�ͽ��ͽ|GνE�ν�ν��ν4�ν��ν�Bν��ͽF�ͽe1ͽ��̽&�̽�̽nt̽P   P   �!̽P̽��̽Q$ͽ�ͽVν��ν�uϽ��Ͻlн�
нm�Ͻ�pϽ��ν{Oν�ͽͽ(�̽�L̽� ̽P   P   ��ʽ�ʽ�>˽�̽�ͽd*ν�RϽ dн&Aѽ��ѽ� ҽ��ѽ�;ѽs\н�IϽ� νh�̽8�˽d9˽�ʽP   P   �ʽ��ʽ6,˽��˽|$ͽt�νi�Ͻ�kѽE�ҽZ�ӽzԽ�Խ�ӽ��ҽ;bѽ��Ͻqzν�ͽ��˽�'˽P   P   d9˽��ʽe<˽��˽�.ͽG�ν�kн.ҽ~�ӽWս��ս�;ֽ��ս$սD�ӽ�#ҽ�aнǪν�&ͽ��˽P   P   8�˽;l˽�m˽�̽�"ͽ�νW�нՔҽB�Խ�:ֽ�y׽"ؽz ؽ�t׽E3ֽ�Խy�ҽ+�нǪν�ͽP   P   h�̽�̽�˽�̽�ͽ-�ν kнL�ҽ��Խ��ֽ7xؽ,�ٽ��ٽ!�ٽJrؽ~�ֽ/�Խy�ҽ�aнqzνP   P   � νK�̽&̽u'̽W�̽='ν��Ͻ6-ҽ~�Խ��ֽ��ؽSIڽ�۽�۽�Dڽ��ؽ~�ֽ�Խ�#ҽ��ϽP   P   �IϽ��ͽ�̽lF̽h�̽,�ͽ}PϽ*jѽo�ӽ;ֽ�yؽ�Iڽ4w۽��۽�t۽�DڽJrؽE3ֽD�ӽ;bѽP   P   s\нsxν�ͽ�k̽
m̽�"ͽ[}ν�bнӨҽ�ս�{׽=�ٽX۽,�۽��۽�۽!�ٽ�t׽$ս��ҽP   P   �;ѽ�.Ͻ6�ͽb�̽L=̽�̽��ͽ�3ϽAѽw�ӽ(�սV%ؽL�ٽX۽4w۽�۽��ٽz ؽ��ս�ӽP   P   ��ѽD�Ͻ�ͽ��̽U̽�̽��̽��ͽ�ϽE�ѽ;Խ�?ֽV%ؽ=�ٽ�IڽSIڽ,�ٽ"ؽ�;ֽ�ԽP   P   � ҽI нy;νN�̽��˽D�˽��˽ �̽�=ν�н�ҽ;Խ(�ս�{׽�yؽ��ؽ7xؽ�y׽��սzԽP   P   ��ѽ@нeRν��̽ �˽�f˽g˽C�˽V�̽�Sν�нE�ѽw�ӽ�ս;ֽ��ֽ��ֽ�:ֽWսZ�ӽP   P   &Aѽg�Ͻ >ν��̽��˽A˽�˽
A˽�˽V�̽�=ν�ϽAѽӨҽo�ӽ~�Խ��ԽB�Խ~�ӽE�ҽP   P    dн�5Ͻ��ͽ\�̽��˽�A˽��ʽ>�ʽ
A˽C�˽ �̽��ͽ�3Ͻ�bн*jѽ6-ҽL�ҽՔҽ.ҽ�kѽP   P   �RϽ��νY�ͽ��̽?�˽i˽	˽��ʽ�˽g˽��˽��̽��ͽ[}ν}PϽ��Ͻ kнW�н�kнi�ϽP   P   d*ν�ͽ4'ͽ��̽̽ �˽i˽�A˽A˽�f˽D�˽�̽�̽�"ͽ,�ͽ='ν-�ν�νG�νt�νP   P   �ͽ��̽��̽�r̽BB̽̽?�˽��˽��˽ �˽��˽U̽L=̽
m̽h�̽W�̽�ͽ�"ͽ�.ͽ|$ͽP   P   �̽�̽�-̽M̽�r̽��̽��̽\�̽��̽��̽N�̽��̽b�̽�k̽lF̽u'̽�̽�̽��˽��˽P   P   �>˽Er˽��˽�-̽��̽4'ͽY�ͽ��ͽ >νeRνz;ν�ͽ6�ͽ�ͽ�̽&̽�˽�m˽e<˽6,˽P   P   �ʽ��ʽEr˽�̽��̽�ͽ��ν�5Ͻg�Ͻ@нI нD�Ͻ�.Ͻsxν��ͽK�̽�̽;l˽��ʽ��ʽP   P   �ȽP�Ƚ�ɽ>�ʽ]�˽Xtͽ~Ͻ�wн�ѽhҽ��ҽ�cҽW�ѽimнq�ν�gͽ��˽��ʽ�ɽ��ȽP   P   ��Ƚ��Ƚ�uɽO�ʽ4̽=�ͽ��Ͻ��ѽޏӽv�Խ�xսsvս6�Խ�ӽ��ѽ��Ͻ�ͽ�̽i�ʽpɽP   P   �ɽ71ɽ؊ɽ/�ʽ�$̽�0ν9�нe�ҽ�ս8�ֽ�ؽswؽ}ؽ��ֽ�ս��ҽ�vн$ν ̽i�ʽP   P   ��ʽ��ɽ��ɽi�ʽ�̽0ν˹нYvӽW!ֽ�uؽ�/ڽ�۽]۽2)ڽ�kؽ�ֽthӽ�н$ν�̽P   P   ��˽ڠʽ�2ʽФʽp�˽��ͽ�н�uӽ�|ֽ�JٽJ�۽ݽ��ݽ�ݽ��۽?ٽ�oֽthӽ�vн�ͽP   P   �gͽզ˽q�ʽP�ʽ<�˽_pͽ��Ͻs�ҽ�!ֽ�JٽRܽ�޽	-߽�*߽�޽�ܽ?ٽ�ֽ��ҽ��ϽP   P   q�ν6�̽`˽��ʽ�c˽��̽uϽ��ѽ�ս�vؽڒ۽�޽�߽�O�A�߽�޽��۽�kؽ�ս��ѽP   P   imн��ͽb̽�˽'˽�̽x�ͽ�uн��ӽ��ֽ�2ڽ�ݽ�/߽�Q��O��*߽�ݽ2)ڽ��ֽ�ӽP   P   W�ѽ��ν��̽^R˽i�ʽ�T˽�̽Y�νѤѽm�Խ$ؽ^۽�ݽ�/߽�߽	-߽��ݽ]۽}ؽ6�ԽP   P   �cҽލϽ�4ͽ׈˽իʽƬʽk�˽�8ͽX�Ͻjҽ�|սT}ؽ^۽�ݽ�޽�޽ݽ�۽swؽsvսP   P   ��ҽ��Ͻ��ͽ�˽T�ʽ�"ʽk�ʽ��˽��ͽ_�Ͻ��ҽ�|ս$ؽ�2ڽڒ۽RܽJ�۽�/ڽ�ؽ�xսP   P   hҽ7�Ͻ�ͽ��˽`vʽ��ɽ��ɽ2wʽ��˽Ӱͽ_�Ͻjҽm�Խ��ֽ�vؽ�Jٽ�Jٽ�uؽ8�ֽv�ԽP   P   �ѽ-�Ͻ��ͽ�˽�pʽ\�ɽ�Hɽh�ɽ�pʽ��˽��ͽX�ϽѤѽ��ӽ�ս�!ֽ�|ֽW!ֽ�սޏӽP   P   �wн �ν�:ͽ �˽gxʽx�ɽɽ�ɽh�ɽ2wʽ��˽�8ͽY�ν�uн��ѽs�ҽ�uӽYvӽe�ҽ��ѽP   P   ~Ͻ��ͽ�̽�˽ɍʽ��ɽ�Iɽɽ�Hɽ��ɽk�ʽk�˽�̽x�ͽuϽ��Ͻ�н˹н9�н��ϽP   P   Xtͽo�̽�̽3Z˽��ʽ�&ʽ��ɽx�ɽ\�ɽ��ɽ�"ʽƬʽ�T˽�̽��̽_pͽ��ͽ0ν�0ν=�ͽP   P   ]�˽��˽Qj˽:"˽i�ʽ��ʽɍʽgxʽ�pʽ`vʽT�ʽիʽi�ʽ(˽�c˽<�˽p�˽�̽�$̽4̽P   P   >�ʽ�ʽ��ʽ�ʽ:"˽3Z˽�˽ �˽�˽��˽�˽׈˽^R˽�˽��ʽP�ʽФʽi�ʽ/�ʽO�ʽP   P   �ɽr�ɽ�:ʽ��ʽQj˽�̽�̽�:ͽ��ͽ�ͽ��ͽ�4ͽ��̽b̽`˽q�ʽ�2ʽ��ɽ؊ɽ�uɽP   P   P�Ƚ�5ɽr�ɽ�ʽ��˽o�̽��ͽ �ν-�Ͻ7�Ͻ��ϽލϽ��ν��ͽ6�̽զ˽ڠʽ��ɽ71ɽ��ȽP   P   2!ƽhnƽqMǽ��Ƚ�tʽ[~̽y�νÒн�,ҽ�7ӽْӽ�2ӽQ"ҽ�н��νEn̽"eʽ	�Ƚ	Dǽ�iƽP   P   �iƽlƽ
/ǽ��Ƚ��ʽ(ͽ��Ͻ4zҽ��Խ�ֽ(j׽Eg׽�xֽ��Խjҽd�Ͻ ͽϟʽ�Ƚu'ǽP   P   	Dǽ��ƽqIǽO�Ƚt�ʽρͽ��нt�ӽ(�ֽLdٽ� ۽�۽��ڽ�Xٽ��ֽ��ӽD�н�pͽ��ʽ�ȽP   P   	�Ƚ��ǽ}�ǽΧȽ��ʽ��ͽ1�н`�ԽTؽ�۽��ݽ�5߽�2߽��ݽ~۽�Bؽ��Խ��н�pͽϟʽP   P   "eʽ��Ƚ�$Ƚ��Ƚ�oʽw%ͽn�н�Խ��ؽ��ܽ3�߽���ʧ�L��b�߽=�ܽ�ؽ��ԽD�н ͽP   P   En̽ʽ��Ƚb�Ƚ*ʽ�y̽[�Ͻ��ӽoTؽg�ܽ<�཭h�u�����:`�}�=�ܽ�Bؽ��ӽd�ϽP   P   ��ν�˽ӱɽ�ɽ��ɽ�˽�ν(yҽT�ֽ��۽�߽gj㽴��F����:`�b�߽~۽��ֽjҽP   P   �н�ͽ˗ʽAUɽWɽ��ʽͽǐн��Խ�fٽ��ݽ���y��e��F�����L�ί�ݽ�Xٽ��ԽP   P   Q"ҽ \ν�s˽��ɽrɽ��ɽz˽eν�,ҽR�ֽ�۽U<߽(��y�佴��u��ʧ⽂2߽��ڽ�xֽP   P   �2ӽ�WϽ�+̽��ɽ��Ƚ7�Ƚ~�ɽ�1̽�_ϽW;ӽp׽l�۽U<߽���gj㽭h�����5߽�۽Eg׽P   P   ْӽ5�Ͻ|�̽�)ʽ�Ƚ�Ƚ��Ƚ`-ʽ�̽��Ͻɘӽp׽�۽��ݽ�߽<��3�߽��ݽ� ۽(j׽P   P   �7ӽ��Ͻm�̽`LʽȽ�ǽW�ǽD�ȽwNʽd�̽��ϽW;ӽR�ֽ�fٽ��۽g�ܽ��ܽ�۽Ldٽ�ֽP   P   �,ҽ�^Ͻ��̽�Mʽ�|Ƚ�Wǽ�ƽXǽ�|ȽwNʽ�̽�_Ͻ�,ҽ��ԽT�ֽoTؽ��ؽTؽ(�ֽ��ԽP   P   н�fνB3̽/ʽ��Ƚ8Yǽ��ƽz�ƽXǽD�Ƚ`-ʽ�1̽eνǐн(yҽ��ӽ�Խ`�Խt�ӽ3zҽP   P   y�ν�ͽ�~˽��ɽn�Ƚљǽ��ƽ��ƽ�ƽW�ǽ��Ƚ~�ɽz˽ͽ�ν[�Ͻn�н0�н��н��ϽP   P   [~̽Ğ˽�ʽ��ɽ��Ƚ�Ƚљǽ8Yǽ�Wǽ�ǽ�Ƚ7�Ƚ��ɽ��ʽ�˽�y̽w%ͽ��ͽρͽ(ͽP   P   �tʽ
 ʽ��ɽ�_ɽpɽ��Ƚn�Ƚ��Ƚ�|ȽȽ�Ƚ��ȽsɽWɽ��ɽ*ʽ�oʽ��ʽt�ʽ��ʽP   P   ��Ƚ�Ƚ��Ƚ�ɽ�_ɽ��ɽ��ɽ/ʽ�Mʽ`Lʽ�)ʽ��ɽ��ɽAUɽ�ɽb�Ƚ��ȽΧȽO�Ƚ��ȽP   P   qMǽ��ǽ�.Ƚ��Ƚ��ɽ�ʽ�~˽B3̽��̽m�̽|�̽�+̽�s˽˗ʽԱɽ��Ƚ�$Ƚ}�ǽqIǽ
/ǽP   P   hnƽ��ƽ��ǽ�Ƚ
 ʽĞ˽�ͽ�fν�^Ͻ��Ͻ5�Ͻ�WϽ \ν�ͽ�˽ʽ��Ƚ��ǽ��ƽlƽP   P   �½b,ý�PĽ� ƽ}ȽU5˽�ν��н@�ҽRԽ�ԽBKԽ��ҽ'�н�ͽ{ ˽�hȽ9ƽ�DĽM&ýP   P   M&ý�)ý-)Ľ�ƽ��ȽF̽�Ͻ�Mӽwֽ��ؽ�ڽ�ڽ��ؽfֽ�8ӽ��Ͻ�̽�Ƚ�ƽ�ĽP   P   �DĽ(�ý�KĽ�ƽ��ȽO�̽��н�@ս:hٽ=�ܽ߽5�߽�߽I�ܽ�Rٽ�(ս��н�̽q�Ƚ�ƽP   P   9ƽ��Ľ�Ľ�ƽp�Ƚ��̽7ѽLֽ	X۽��߽�&�g����^㽳�߽a@۽�2ֽhѽ�̽�ȽP   P   �hȽ�(ƽOgŽ�/ƽ�vȽ�̽-�н�Kֽrܽ�j�-��I�����U�软��HU�e�۽�2ֽ��н�̽P   P   { ˽$�ǽ�UƽrYƽ��ǽ0˽��Ͻ@սnX۽�k�h��!��c	����н�HU�a@۽�(ս��ϽP   P   �ͽ��ɽ�rǽB�ƽ�xǽ��ɽ�ν�Lӽ3iٽh�߽��彩��6-R��$�꽯�彳�߽�Rٽ�8ӽP   P   '�н`�˽�Ƚ0�ƽ��ƽ��Ƚ��˽��н�xֽ��ܽ�,�+��!�UｵRｓ�U��^�I�ܽfֽP   P   ��ҽ/�ͽ��ɽ�^ǽыƽ�cǽw�ɽ[�ͽ��ҽ��ؽ�߽��低��!�6-�c	�����佹߽��ؽP   P   BKԽMϽW�ʽ��ǽ/<ƽ�=ƽ��ǽ��ʽ�Ͻ^WԽ1ڽ��߽���+�轩��!��I��g��5�߽�ڽP   P   �Խ��Ͻoo˽%Ƚ�ƽ6UŽCƽ�!Ƚv˽�Ͻ��Խ1ڽ�߽�,����h��,�彞&�߽�ڽP   P   RԽ9�Ͻ;�˽NȽ��Žh�Ľ�Ľ�ŽAQȽ��˽�Ͻ^WԽ��ؽ��ܽh�߽�k��jὩ�߽=�ܽ��ؽP   P   @�ҽ�Ͻ�t˽+PȽr�ŽeĽ�ýgeĽW�ŽAQȽv˽�Ͻ��ҽ�xֽ3iٽnX۽rܽ	X۽:hٽwֽP   P   ��н��ͽT�ʽ�#Ƚ��ŽYfĽl�ýs�ýgeĽ�Ž�!Ƚ��ʽ[�ͽ��н�Lӽ@ս�KֽLֽ�@ս�MӽP   P   �νH̽��ɽ��ǽ,ƽθĽ��ýl�ý�ý�ĽCƽ��ǽw�ɽ��˽�ν��Ͻ-�н7ѽ��н�ϽP   P   T5˽�ʽ��Ƚ
kǽ�Dƽ:[ŽθĽYfĽeĽh�Ľ6UŽ�=ƽ�cǽ��Ƚ��ɽ0˽�̽��̽O�̽F̽P   P   }ȽqȽ��ǽ~ǽ��ƽ�Dƽ,ƽ��Žr�Ž��Ž�ƽ/<ƽыƽ��ƽ�xǽ��ǽ�vȽo�Ƚ��Ƚ��ȽP   P   � ƽ�8ƽeƽ��ƽ~ǽ
kǽ��ǽ�#Ƚ+PȽNȽ%Ƚ��ǽ�^ǽ0�ƽB�ƽrYƽ�/ƽ�ƽ�ƽ�ƽP   P   �PĽ�ĽmtŽeƽ��ǽ��Ƚ��ɽU�ʽ�t˽;�˽oo˽W�ʽ��ɽ�Ƚ�rǽ�UƽOgŽ�Ľ�KĽ-)ĽP   P   b,ý�ý�Ľ�8ƽqȽ�ʽH̽��ͽ�Ͻ9�Ͻ��ϽMϽ0�ͽa�˽��ɽ$�ǽ�(ƽ��Ľ(�ý�)ýP   P   6d��
辽d��e�½��Ž�zɽ�Fͽ��нi�ӽP�ս�|ֽ$�ս��ӽ��н2,ͽ�_ɽ��Ž\�½�T��:྽P   P   :྽�侽2��c�½�Kƽ��ʽ��Ͻ�iԽ��ؽ��۽	�ݽe�ݽ��۽��ؽ�MԽ�oϽN�ʽ*2ƽ]�½�%��P   P   �T�������]��д½sƽ�Z˽�ѽ�׽��ܽ�����c�彀��p��ܽw�ֽ��н�<˽3Zƽ]�½P   P   \�½=�������H�½Hƽ�Y˽�ѽ��ؽ�|߽���Rk��������Y�K��N\߽tdؽxѽ�<˽*2ƽP   P   ��Ž��½���*�½�Ž֭ʽ7ѽ��ؽ.o���Eq����/e�.�B���L�tdؽ��нN�ʽP   P   �_ɽ�&Ž� ý�ý�3Ž�tɽ��ϽW׽`}߽���'�ｓl��s��������[����B��N\߽w�ֽ�oϽP   P   2,ͽX�ǽ�wĽ�Zý�Ľ��ǽ�BͽiԽ�ܽ���OI��o���4��6���b)���[��.�J���ܽ�MԽP   P   ��н�tʽ.ƽ�ý��ý�ƽ��ʽ��нV�ؽ$�ὒs�Cz�~�������6�������/e��Y�pὕ�ؽP   P   ��ӽ-�̽��ǽ�^Ľ�Hý�dĽ��ǽ��̽U�ӽ�ܽ��U ���~����4��s��������콀�佇�۽P   P   $�ս۩νf�ȽL�Ľ,�½e�½\�Ľ��Ƚa�ν6�ս�ݽ	��U �Cz��o���l���q����c��e�ݽP   P   �|ֽe�Ͻ�ɽ�dŽt�½ڹ��I�½kŽ��ɽ��Ͻ��ֽ�ݽ�佒s�OI�'��E�Rk���	�ݽP   P   O�սi�Ͻ�#ʽۨŽˇ½��������Պ½��Ž�)ʽ��Ͻ5�ս�ܽ$�Ὅ�彉���罗�彯�ὺ�۽P   P   i�ӽ˵ν��ɽ��Ž�~½����ۿ�v�����½��Ž��ɽa�νU�ӽV�ؽ�ܽ`}߽.oཛ|߽��ܽ��ؽP   P   ��н��̽B�ȽwlŽ6�½I�����������v���Պ½kŽ��Ƚ��̽��нiԽW׽��ؽ��ؽ�׽�iԽP   P   �Fͽ�ʽ�ǽ��Ľx�½�����ݿ������ۿ�����I�½\�Ľ��ǽ��ʽ�Bͽ��Ͻ7ѽ�ѽ�ѽ��ϽP   P   �zɽ��ǽ/#ƽ�mĽ��½��������I����������۹��e�½�dĽ�ƽ��ǽ�tɽ֭ʽ�Y˽�Z˽��ʽP   P   ��Žp>ŽËĽ��ý�Uý��½x�½6�½�~½ˇ½t�½-�½�Hý��ý�Ľ�3Ž�ŽHƽsƽ�KƽP   P   e�½F�½�ý�ký��ý�mĽ��ĽwlŽ��ŽۨŽ�dŽL�Ľ�^Ľ�ý�Zý�ý*�½H�½д½c�½P   P   d�����U����ýËĽ/#ƽ�ǽC�Ƚ��ɽ�#ʽ�ɽf�Ƚ��ǽ.ƽ�wĽ� ý��������]��2��P   P   
辽򙿽���F�½p>Ž��ǽ�ʽ��̽˵νi�Ͻe�Ͻ۩ν-�̽�tʽX�ǽ�&Ž��½=��������侽P   P   �����]���E���W��&g½�*ǽ�:̽�ѽ�ս��׽H�ؽ��׽�սh�н̽#ǽ�F½�<���2���S��P   P   �S��`Y������L��1�½�Ƚ<NϽX�ս�۽hJཻ�⽅�⽭5ཽ�۽7�ս�%Ͻp�Ƚ��½�2������P   P   �2��[4���>��eI���0ý�ɽ3\ѽ��ٽuj�;轉h����X���罌C��^ٽ�0ѽX�ɽ�ý�2��P   P   �<��滽컽�N����½_�ɽ�ҽz�۽�,彮����;��t2��W������A ��W۽F�ѽX�ɽ��½P   P   �F½�[��x��h��V^½c�ȽlZѽw�۽��!� ��T �$�� �� ������O��W۽�0ѽp�ȽP   P   #ǽ�p��|���M������g#ǽ�JϽ��ٽ].�$�%���A�R����A5�/������A ��^ٽ�%ϽP   P   ̽��ĽV������c���L Ž�6̽��ս�m�_���&���C����������A5�� �����C�7�սP   P   h�н/uȽ�½��������d�½u�ȽSѽ��۽�
轌���� �"��	������� �V�����罽�۽P   P   �ս��˽v�Ľ�h�������p����Ľ��˽'!ս�T�Qx콣N���.�!�����R��$�s2���X콭5�P   P   �׽�ν�rƽj-��E���z���<7��k�ƽT0ν��׽l�⽤N��� ��C��A�T �;������P   P   H�ؽ`rϽ��ǽw����8�����o=������*�ǽx�Ͻ�ؽl��Qx콌����&��%��� �����h콺��P   P   ��׽�wϽ�Ƚ,½�����a�����B3½�Ƚx�Ͻ��׽�T��
�_��$��!���:�hJ�P   P   �ս_+νN�ǽ�/½���񂻽����5���S��B3½*�ǽT0ν&!ս��۽�m�].���,�uj��۽P   P   �ѽ�˽w�ƽ\���L������1���0��5����������k�ƽ��˽Sѽ��ս��ٽw�۽y�۽��ٽX�սP   P   �:̽�Ƚ)�Ľ�<��\B��������1������a��o=��<7����Ľu�Ƚ�6̽�JϽlZѽ�ҽ3\ѽ;NϽP   P   �*ǽ�	Ž4�½�{�����x��������񂻽������z����p��d�½L Žg#ǽc�Ƚ^�ɽ�ɽ�ȽP   P   &g½��������d���~
�����\B��L��������8��F�����������c������V^½��½�0ý1�½P   P   �W���u��0���b!��d����{���<��]����/½,½x���k-���h���������M���h���N��eI���L��P   P   �E��I���="��0�������4�½)�Ľw�ƽN�ǽ�Ƚ��ǽ�rƽw�Ľ�½V���|���x��컽�>�����P   P   �]��)A��I����u�������	Ž�Ƚ�˽`+ν�wϽ`rϽ�ν��˽0uȽ��Ľ�p���[��滽[4��`Y��P   P   ej���>�����}���xӽ�Ľ?�ʽ ?ѽ��ֽ�cڽX�۽	Sڽ%�ֽkѽ��ʽ�ýN����t��[���H2��P   P   H2���8���]��a���(����?ƽ6�ν0�׽=�߽��iy�p�7�归�߽>�׽�ν�ƽ�t��tm��6I��P   P   [���nK��^��������澽�rǽn�ѽr�ܽ)�����)���X��Q��Z��pv��ܽ�tѽ�>ǽK���tm��P   P   �t��+o��*w������Ě���pǽ��ҽÍ߽����T��z�����h�� �����N߽�oҽ�>ǽ�t��P   P   N��������ⶽ����`ɽ�	:ƽ֬ѽߍ߽�������>����	���]�	�Lj������N߽�tѽ�ƽP   P   �ýr���߸��渽����~Ľ!�ν#�ܽ
���������1�Ң�W��P�n���������ܽ�νP   P   ��ʽ��SS��)k���a���/����ʽ�׽���:]�����4�My��W��m�P�Lj�� ��pv�>�׽P   P   kѽ�Ž��^7��:>��:#��z�Ž@ѽN�߽�𽌂�w�	�M��*]��W�V��]�	��h�Z�𽑵߽P   P   %�ֽfʽ�����6���[���A������� ʽ��ֽ�(��?��Z*�k��M��My�Ң�����Q��7��P   P   	SڽwKͽY#ýE?���Ǹ�\̸��L��A8ý�gͽtڽ��iz��Z*�v�	��4��1���	���X��p�P   P   W�۽�Ͻ��Ľ���(w��B춽}���(����Ľ�0ϽE�۽���?����������>��z�~)��hy�P   P   �cڽ� ϽRQŽf����T������ۭ��+[��ǥ���^Ž�0Ͻtڽ�(���:]����������T������P   P   ��ֽ3_ͽ��Ľџ���O��������'���S��ǥ����Ľ�gͽ��ֽM�߽���	��������(��<�߽P   P   �>ѽ ʽ!8ý(���Z�����g���g��'��+[���(��A8ý� ʽ@ѽ�׽"�ܽލ߽Í߽r�ܽ0�׽P   P   ?�ʽ)�Ž
���2R���������������g������ۭ���}���L������z�Ž��ʽ �ν֬ѽ��ҽn�ѽ5�νP   P   Ľ.:��k/���N���׸�F���������������C춽\̸��A��:#���/��~Ľ:ƽ�pǽ�rǽ�?ƽP   P   xӽ�-���s���P���m���׸������Z���O���T��(w���Ǹ��[��:>���a������`ɽ�Ě���澽'���P   P   }���w���4��������P���N��2R��(��џ��g������F?���6��_7��)k���渽������������a���P   P   ���t�������4���s��k/�����!8ý��ĽRQŽ��ĽY#ý������SS��߸��ⶽ*w��^����]��P   P   �>��1[��t���x���.���/:��)�Ž ʽ4_ͽ� Ͻ�ϽxKͽgʽ�Ž��s�������+o��nK���8��P   P   �&��.��_2��u!���ͷ��ۿ�)�Ƚ"Oѽ��ؽʰݽ�o߽C�ݽJ�ؽ ѽ�mȽĠ��֙�����������P   P   ���['���ի����޸�^�½�0ν� ڽ�7彬���򽠋�������ٽ��ͽ��½s�������߻��P   P   ���dy���'������?��
_Ľ�ѽ3�\� '��]�$������������c��O�ѽ@Ľ;
������P   P   ����!���+������ظ�	]Ľ�Gӽ ����������/��,��Ύ��|��3��z�S�ҽ@Ľs���P   P   ֙������ꮽd%��6·�W�½��ѽ[�但3�����{X����F����#������z�O�ѽ��½P   P   à��h���f���p���;��$ҿ��-ν��ٍ��=�����L�џ"��"�J1�Ħ�#���3��c����ͽP   P   �mȽ��������ݘ��+���Ƚ�#ڽ��ҧ���bQ��~%��n(�hm%�J1�����|�����ٽP   P    ѽ�½x������$���'���5½mRѽZB�y:��X���f���"�>w(��n(��"�F�Ύ��������P   P   I�ؽ�ǽ񞻽m�����j{�������ǽA�ؽ7����������"��~%�џ"����,�������P   P   B�ݽm̽Ҷ��ϵ��b���h���ൽ=Ӿ��7̽��ݽ��M�����f�bQ��L�zX�.��#�����P   P   �o߽�|ν:���%�����R�������������ν��߽���X�����������]����P   P   ɰݽ�ν�������������*�������0��������ν��ݽ7��y:��ҧ�=����� '�����P   P   ��ؽ�*̽%���-������ެ�O���⬽����0��������7̽A�ؽYB彯�؍���3�����[�7�P   P   !OѽW�ǽ�о�V	�����ᬽ�Ѫ��Ѫ�⬽�������=Ӿ��ǽmRѽ�#ڽ��Z�����3�� ڽP   P   (�Ƚ�:½����浽��젭�K����Ѫ�O���*�������ൽ�����5½�Ƚ�-ν��ѽ�Gӽ�ѽ�0νP   P   �ۿ��$��(5�������u��T%��젭�ᬽ�ެ����R���h��j{���'��+��#ҿ�V�½]Ľ	_Ľ]�½P   P   �ͷ�bL��?���7:��R#���u��������������b������$��ݘ���;��6·��ظ��?���޸�P   P   u!��t9��:����2��7:������浽W	��-�������%���ϵ�m���������p��d%��������
��P   P   _2���@�����:���@���)5�������о�&�������;���Ҷ��񞻽y������f���ꮽ�+���'���ի�P   P   .�������@��u9��bL���$���:½X�ǽ�*̽�ν�|νn̽�ǽ�½��h������!��dy��['��P   P   �����Ý��r������毽�*����Žѽ��ڽr�Ὕ&�ۧ���ڽ��н2NŽ,๽#���(U��{N�����P   P   ��������K����L�������̽��ܽ2콇��/���]�������B��،ܽǎ̽��������]���栽P   P   {N��S���e��h����α������ѽ�R��?�����o�����X�#����������ѽ����ɉ���]��P   P   (U��b������S{��tE��_��Ӿӽ?���� ��:�# �� �����>��뽡Uӽ�������P   P   #����g����������ٯ�j���ѽe�뽋������W#�E�-�0�1��-��%#�ą������ѽ����P   P   ,๽@����ŧ��ҧ�eޭ�� ����̽�U潈��'���&�o�5�7)>��>��n5�.s&�ą�=�����Ǝ̽P   P   1NŽ#��D���c����ǫ��S��8�Ž7�ܽ�L��!��	b#���5���B�ݨG��B��n5��%#�������،ܽP   P   ��н�����-���쩽�����O���4��ѽN#콱��<L���-�=>���G�ݨG��>��-���"��A��P   P   ��ڽ^ĽZĴ����c���긫�&괽̕Ľd۽�=������A �v�1�=>���B�6)>�0�1�� ��X�����P   P   ڧ�.*ʽ�̸�o{���什�����������]ʽd���������A ���-���5�n�5�E�-�# ����\���P   P   �&��bͽ���D	������3������p ������x�ͽ�W�������<L�	b#��&��W#� :�o�.���P   P   q��unͽ���������q��v��+������뵼�w�ͽd���=�����!��&����� ��������P   P   ��ڽKKʽ��������L���j���u������g�����������]ʽc۽N#콃L�����������?��1�P   P   ѽ��Ľ�츽q������㝢�A!���!�����,���p ����̕Ľѽ7�ܽ�U�d��>�뽑R���ܽP   P   ��Ž�8���@������ny�����A!��u���v����������&괽�4��8�Ž��̽��ѽҾӽ��ѽ�̽P   P   �*��`��X]���ǫ����~>��ny��㝢�k����q���3������긫��O���S��� ��i�^���������P   P   �毽�𭽞ޫ����lŨ�����������L����������什c��������ǫ�eޭ�ٯ�sE���α��L��P   P   ���蘧���X�������ǫ�A���r�������E	��p{������쩽c����ҧ�����R{��h���K���P   P   �r��k���`ۤ��𧽟ޫ�Y]����츽������������̸�[Ĵ��-��E����ŧ���������e����P   P   �Ý�Ij��k���蘧���`���8����ĽLKʽvnͽ�bͽ/*ʽ^Ľ����#��@����g��b���S�����P   P   ������-��L�������n�����lн�]ݽ�����齲p潼ݽ��Ͻ�������B��}���Ǔ�#y��P   P   #y�������u��Ta���^��Q��E�ʽ��߽���������v�����G��x߽�.ʽy綽����!��&O��P   P   �Ǔ��f��n䓽�[���������Oѽy��H���a����,n�����(�ȴ�63콁�нU��������!��P   P   }���<���L��D=��IW���
���ӽ�����;q��Z/�9�8�;z8�I#/�,$�;�@a�E)ӽU������P   P   �B�����L̗�E4������EK��OѽO���S�5�&���=��ON�JyT�0#N�#M=�w�&����@a��нy綽P   P   ���rѢ��{��-������3e����ʽ��S��� '���B��2[� �i�V�i�S�Z���B�w�&�;�63콽.ʽP   P   ������ZJ��9����i��%Q�����j�߽^��~�C�=��>[�n�q���y�\hq�S�Z�#M=�,$�Ǵ�x߽P   P   ��Ͻ���w꥽Z,��3:������U��"н����u��u/�ZpN�1�i��z���y�U�i�/#N�H#/��(��G��P   P   �ݽ^���Q���Kd��P����|��T��ۿ��xݽ������8���T�1�i�n�q� �i�IyT�:z8�������P   P   �p潭'ǽl簽Iɢ��������.碽���?lǽ���b������8�ZpN��>[��2[��ON�9�8�+n��v�P   P   ��齦g˽݀���֤��Ǜ��ؘ�,כ����������˽��b�����u/�C�=���B���=��Z/�������P   P   ����v˽�ӵ�K	���ӛ��ܖ�a▽D䛽�#��'����˽������u��~�� '�4�&�:q��a���P   P   �]ݽ&Rǽ7�������䛽���������񛽳#������?lǽ�xݽ����^�S���S����H�����P   P   kн�п�����줽�ݛ��𕽧���	������D䛽��������ۿ�"нi�߽��N����x�콱�߽P   P   ���iW���﫽ꢽ�ٛ��䖽�����������b▽,כ�.碽T��U�������ʽOѽ�ӽ�OѽC�ʽP   P   �n���]��g#��+�������䘽�䖽���ܖ��ؘ�����|�����%Q��2e��DK���
�����Q��P   P   ������{����U��Nٜ�����ٛ��ݛ��䛽�ӛ��Ǜ�����P���3:���i���������HW������^��P   P   �L��N��ϭ������U��+���ꢽ�줽���L	���֤�Jɢ�Ld��[,��9���-���E4��C=���[��Ta��P   P   ,󓽉h������Э��{���h#���﫽���8����ӵ�ހ��m簽R���w꥽[J���{��L̗��L��n䓽�u��P   P   �������h��N�����]��jW���п�(Rǽ�v˽�g˽�'ǽ_���������rѢ�����<���f������P   P   ��x��F|�h9���݋�)������m{����ͽ��߽��ȅ���t:߽v~ͽ
������UǗ���������|�P   P   �|��2|�@���j ��g�����a�ƽ��⽈;��`i��,�,��6�����O⽄7ƽۙ������^���x��P   P   ����>��P)��b����7������ �Ͻ\P������!��/0��l5�l 0���!�#�y���ν���͚�^���P   P   ����寄�NÄ�c̋�\_������ҴҽG���f��k5��
N�~�\��\�#�M��4����l����ѽ������P   P   UǗ�����G����������^���ϽaJ���m���@���d��L�����,(���cd�2p@�����l����νڙ��P   P   ����I̔�	���C���	�����ƽ�X��Jm�� A���m��X��������^!��b�l�2p@���y��7ƽP   P   	��I���ő��<��푽rh��v|����⽕���~5���d��b��O������&��^!���cd��4�#�O�P   P   t~ͽ{���N���HV���g��Dܘ��ν�\���"��2N��f��].�����������,(��"�M���!�����P   P   r:߽����䟽O)���̍�:H��C#��.��"�߽���`0�A�\�񸅾].��O��������\�k 0��6�P   P   ���·½.k��]:������+��E`��d���j�½\M��]���5�A�\��f���b���X���L��}�\��l5�+�P   P   Ņ�Ƚ����ޗ�Y��0���-��h���>���eȽ���]�`0��2N���d���m���d��
N��/0��,�P   P   ��C-Ƚ�����i���Q��������Rg��ˌ���䬽�eȽ[M콄���"��~5�� A���@��k5���!�^i�P   P   ��߽��½s���r��t�������U��홆�����ˌ���>��j�½!�߽�\�����Im��m��f����;��P   P   ��ͽ���E��������\��=��� J��yL��홆�Sg��h��d���.���ν��⽸X��_J��G��ZP�����P   P   l{��Q쬽|"���_���,��C���[V�� J���U�����-��E`��B#��u|����ƽ�Ͻдҽ��Ͻ_�ƽP   P   �����s��:阽fU���8������C���>����������1����+��:H��Dܘ�qh���]�������������P   P   )�������Q���ꍽ�8���,���\��t���Q��Z������̍��g��푽�	�����[_���7��g��P   P   �݋�΋�b8��*h��Q���fU���_�������r���i���ޗ�^:��P)��HV���<��C������b̋�b���i ��P   P   g9���ℽ4ԇ�b8��	��;阽}"��G���t�� ������/k���䟽O����ő�	���G���NÄ�O)��@���P   P   �F|��]���ℽ�΋�����s��R쬽�����½E-Ƚ�ȽЇ½���|���J��I̔�����寄��>���2|�P   P    N��HR���]�Wq��
������	��-�ɽ�ཝ��'���GU�+���Oɽ�r���������(�p�Y9]��R�P   P   �R��0R��}\�Ͽq�=�k�������4�!������Fz����J��g�V߿�� ���D��q�Q\�P   P   Y9]�{�V���]���q�����<�����˽�o���W�E6���K�'|S��BK��5����Wm��;�ʽ	K��<B��q�P   P   (�p�F�`��a��1q���+���M�Ͻ ����)��wS���y��Ո������fy���R�B7)��j��Ͻ	K���D��P   P   ���܀p���g���p���������Y�˽"����/�VKe�ۖ��|O���������5���zd���.��j�;�ʽ� ��P   P   �������χq���q�#V��D	��p���K{���)�ZUe�[▾����Ҿ��Ҿ
���^l���zd�A7)�Vm��U߿�P   P   �r����������t��}�����H���F彩h���S������)������X𾅧�
���5����R�����g�P   P   �Oɽ����҇���y���y�u���R��Y�ɽ����j6��%z�wz���Ӿ�|��X���Ҿ����fy��5�J�P   P   )��2��b���Cp����v�W������������*��-�o�K�����簾Ӿ�����Ҿ���������BK����P   P   DU����ʘ��S����u��v�؂��#��>�����$����S����wz���)����{O���Ո�%|S�Dz�P   P   $�����½v���ư���~v�d�n�0�v�Y⇽�ڞ�d(ý���$��o�K��%z�����Z▾ۖ����y���K���P   P   ���k�½e���ը���yw�V�j�}�j��w�wՉ�|�d(ý����-��j6���S�YUe�UKe��wS�E6���P   P   �ཡܻ���������m�w�{�h��c�k�h�'!x�wՉ��ڞ�>���*ὀ���h��)���/���)��W� ��P   P   +�ɽ�s������͇�w�w��h��a�I�a�l�h��w�Y⇽#������Y�ɽ�F�I{��!������o���4�P   P   �	���L��$���W}���v���j��c��a��c�~�j�1�v�؂�������R��G��o���W�˽K�Ͻ��˽|���P   P   �������������v��n���j��h�|�h�X�j�e�n��v�W���u������C	������*���;���i���P   P   �
���j��J���0z��w��v��v�z�w�p�w��yw��~v���u���v���y��}�"V������캉�����;�P   P   Wq�?q�r�.�t��0z�����X}���͇�����֨��Ȱ���S��Dp����y���t���q���p��1q���q�Ϳq�P   P   ��]��Sa���g�r�L����&����������g���x���ʘ�d����҇���Їq���g��a���]��}\�P   P   �HR�5W��Sa�Aq�k������L���s���ܻ�n�½��½���4�������������݀p�F�`�z�V��0R�P   P   ���k� ���,���B�sqc�.���ƣ���½�ཷ��������V��߽����"��ge��slb���A��},�Fv �P   P   Fv �1� ���+�yGC���i�[��f綽DH彪��O�!�Q/�q�.�<m!�,�sD�����M����h�?}B��B+�P   P   �},�F�%���,�#;C�)l��I��\�Ľ`����'��"O�,Rn��?z���m�N}N�L�&��y�ý�w����j�?}B�P   P   ��A�ii0��0�ɔB�/�i�OH���#ʽ͹
�'k=�o>z������I��	!��P����Dy�j�<���	�� ɽ�w����h�P   P   rlb��A�o�7�K'B�Wc�r
��U�ĽW�
���E�r�4�����3'��N��8����$��K�D���	�y�ý�M��P   P   fe��FZ��B��C���Z�� ��[�����w=��Ɋ�ƾ� �$�������JFž�$��j�<�����P   P   !��a�y�ԑR�_�F�@S�,�z��ϣ�`�.�'�mdz�ô��(���*��.<��O*���8����Dy�K�&�rD�P   P   �����?���f�6M�KEM�M�f�ʏ���½~���UO�'���]�_��X<��.<����M��O���M}N�,�P   P   ߽rѡ�I{���U��J��GV��|��d��T�m"���n�>���Я��_����*�#��2'��!����m�:m!�P   P   �V���^��l���Ȭ_�a�J���J�v`�ᇽ�뱽���`\/��z�>����]�(�� ��㾲I���?z�o�.�P   P   ����(`������h�@L�ѸC�|L��h��ٺ�I(��`\/���n�'��´��ƾ3�������*Rn�O/�P   P   ����_}���7���m�N��@��$@�TTN�y�m����ٺ����m"��UO�mdz��Ɋ�q�m>z��"O�M�!�P   P   ��3���m���W0m�F�N��>��9�U�>�cO�y�m���뱽T�~��-�'��w=���E�%k=���'����P   P   ��½C��F���]h�'N�|�>�q7��z7�V�>�UTN��h�ᇽ�d����½`����V�
�̹
�_��AH�P   P   �ƣ�����#�{��`�!hL�Z@��}9�q7��9��$@�|L�v`��|�ʏ��ϣ�Y�S�Ľ�#ʽY�Ľd綽P   P   +����z�V�f�yUV�p�J�C�C�[@�~�>��>��@�ӸC���J��GV�M�f�*�z�� ��p
��MH���I��X��P   P   oqc�=[��0S��zM��J�q�J�#hL�'N�J�N�N�@L�d�J��J�LEM�?S���Z�Wc�,�i�)l���i�P   P   ��B��aB��lC�r�F��zM�{UV��`�]h�\0m��m�h�ˬ_���U�8M�_�F��C�J'B�ǔB� ;C�wGC�P   P   ��,��0��8��lC��0S�Y�f�'�{�I���p����7������n���I{��f�֑R��B�n�7��0���,���+�P   P   k� �p�%��0��aB�@[���z������C��6���c}��+`���^��tѡ��?��c�y�FZ��A�ii0�E�%�0� �P   P   �ǼQ:ϼ��{����/�5pb����j����ڽ}}���i��
����ٽ4���@Ő�}a�
�.���
���R�μP   P   S�μϼ6W�,k��6�w����������,�0>���=��,��9��`߽j���Su�X�5�����V�P   P   �缻Uټ&��X_�Ô9�M�����},�MP4�9�i��䔓�s�����h��b3�:\�E���`����C8����P   P   ��
���ＵI�/��R�6�����;������|Q�ɖ��ݓ���N߾�߾>���;䒾�DP�&��%ݽ�`���W�5�P   P   	�.�ו
�^��/��/�
w�l������z�\��ɧ���>��-�������ᦾI}[�&��D����Su�P   P   za�c�%�#	�I�a�&��lb��$��6��Q��ӧ�����A���u���u��A�����ᦾ�DP�9\�h��P   P   >Ő��I������� @�9�J�!���r���l4�ɰ���"��A�<��4���ދ��A����;䒾�b3��`߽P   P   1����t��14�˚�4��5�4�{Uu�j���}��tj�e���r���dv� f��4����u����<�����h��9�P   P   ��ٽ����)M���#�E2���#��M�P���{�ڽp�,��5��O�߾.��dv�<����u��-��߾r����,�P   P   ������Id�S�/���r��A-0��*e�y2��1�����>�h��O�߾r����A���A��>��N߾┓���=�P   P   �i��%k��� u�J:�����Y�O�:�H�u�(���> ���>��5��e����"�����ۓ���->�P   P   y}������h{�9@�k�)�����f���@��|�(���1���p�,�sj�ɰ���ӧ��ɧ�ǖ��6�i�|�,�P   P   �ڽd袽�pu��P@�CQ � ��]�
����x� ���@�H�u�y2��z�ڽ|���l4��Q�x�\��|Q�KP4����P   P   f����s���d��X:�j+�`��	��)	�����f�P�:��*e�P���i���p��6�������{,����P   P   
���3u�c�M�10��7����N�
�	�^�
���Y�B-0��M�yUu�����$��j����;������P   P   0pb���J���4���#�s�������b��#��,�����t����#�5�4�7�J��lb�
w����J���w�P   P   ��/�ѷ&�	g���a�u���7�m+�GQ �o� ���G2�4�� @�_�&��/�O�6���9��6�P   P   y���K�+��P�����#�50��X:��P@�9@�O:�W�/���#�͚����I�.�-��V_�)k�P   P    ����� �-��g���4�h�M�"�d��pu�h{�� u��Id�.M��14����$	�^���I�#��3W�P   P   P:ϼ�ټ	��K�Է&���J�3u��s��h袽����)k����������t��I�e�%�ؕ
���ＺUټϼP   P   B���k��BS�����`��Q�*���r������ͽ�W�i)�����s�̽�����&q� )�dg�C��Q��Z�P   P   �Z��
�F�N�g������R�@�8���PԽi��л2��H��_H�*2������ҽ}d��u?����	���hlL�P   P   Q��c3�ʿR�6S��N]��w9N�����@ ��4<��!��x8��䨾}ٜ��#�;�v����D��� L�����	���P   P   C���Ta�nEb��������6;N���)��k�`��稾y6���
��
��U�L����f_�n��	`��� L����P   P   ag�'ɗ�@���ژ�n����@���������xo�$�ľ�y��4X��u��W�����þt�m�n���D��s?�P   P   )��NҼ�͛��X��� Լ�*�:��� L �a�j�ľI�*�����������Db��p�)��þ�f_�t���{d��P   P   �&q����ü�k��0$ļ���s��*Խ�V<�i	����*�����e��Db�����K���;���ҽP   P   񹢽��?��z���/��f�������3A�*ڣ���[L������X�Β��2���e������W��U群#����P   P   n�̽�Sq����#ּA����ּ�����r�L�ͽp3����(b��rv�Β��
������u� �
�{ٜ�
*2�P   P   }��=썽�w1�wp� ļ"~ļ����(s2�������n%I��s��(b��X�*������4X���
�䨾�_H�P   P   c)��#r���D�fg�mKϼ���Q�ϼP�źE�������n%I���������H�*��y�v6�v8���H�P   P   �W�O���@�K����*�ؼ#��"\���gټ�Z��L������p3�ZL��h	��i�ľ"�ľ�稾�!��ͻ2�P   P   ��ͽlS��
 E�Z���Zܼ���0糼%x��ݼ�Z�źE�����K�ͽ���V<�a��xo�h�`��4<�f��P   P   ����qr��2�����ؼ��~���vʱ�'x���gټP�(s2���r�(ڣ��*Խ�K ����'���@ �KԽP   P   ��r�A�����#��-�ϼB���������4糼%\��T�ϼ��������3A��s�7������������4���P   P   K�*����/�����ּ gļT���E�������)�����&~ļ��ּ������*���@�1;N�q9N�L�@�P   P   W�漋-Լ3Zļ4�B���#gļ2�ϼ�ؼ�Zܼ4�ؼvKϼ� ļA��i���/$ļ� Լh������E]��w���P   P   z���0;��8ޜ�V��7���ּ�#�����a�����lg��p�+ּ�/���k���X���ژ�����0S���f��P   P   �BS�DRc��Ё�:ޜ�9Zļ8�������2� E�I�K��D��w1�����z���ü�͛�?��iEb�ÿR�>�N�P   P   }k�$�4�HRc�5;���-Լ ��A��qr�qS��T���(r��B썽�Sq���?����NҼ)ɗ��Ta��c3��
�P   P   �_<m��;;�;#+���=���Ҽ��6�p������Yڽ��o�ٽ�4��D��ɻ4�a�ϼ�9�h�.Y�;ε�;P   P   ̵�;{[�;O�;MJ�D�Z������Bk�Y"��}s��V0��wI�L8I��/����Ș����h�R	���GU������;P   P   -Y�;�q�;L�;�
�f�2���������:�����姾���t���t���9����kx��gv�1/`�
���P   P   P���G;�D;]���r�Z�����ʑ�c=��Te�C��	���!��� �N$� �ԕc�C�5��fv�~GU�P   P   �9�V��\�v:	� ���=�� ����@A��Sv���ؾ�5�����0��~%���i4�+׾@Zt�C�jx��M	��P   P   Z�ϼ8�9A)� �-������Ҽ:bk��#��ie���ؾ��M��+���l
�X
����aL�*׾ӕc������h�P   P   û4��y��� ����H��顼:�6�%I���;�a7��ü5��Z����.��v^�N�-�����i4����9�Ř��P   P   @��*����n�S}��w���r����	?��ǟ��J��Z�������
��^��v^�W
�}%��M$��t�����P   P   �4��H-8�˞����;��	��=�|�����9��s��z�0��J��ɣ!��ǜ���
��.��l
�.���� ��t��޳/�P   P   i�ٽf��o����S&�`'�.>�����&h��ڽfJ�����ɣ!�����Z���+�������!���H8I�P   P   ���������4����H��'�:J�K���+������Zw�fJ��J��Z��¼5���M��5����姾�wI�P   P   �Yڽ+��F�������}d�0U1���1��f����fl������ڽy�0��J��`7����ؾ��ؾ@������V0�P   P   ����ig����䰼�6o�z1:�Ki+��;���p����+���&h��s��Ɵ��;��ie��Sv��Te���:�zs�P   P   k���S9���@���-�d�=:�c�*��*��;��f�M�������9�?��#I���#�>A�`=���S"��P   P   ��6����� ��릁��2I��1�! +�h�*�Si+���1�:J�0>��|������7�6�5bk�����ʑ�����Bk�P   P   ��Ҽ�����q�� =���&�c�&��1�I:��1:�?U1��'�k'���=�r��顼��Ҽ� ����,������P   P   ��=�<���u�R��XP	���&��2I�?�d��6o��}d���H��S&��	�����H������=�a�Z�	f�/�Z�P   P   �*�b
�a1�|���`��� =�����M���䰼����	5�����ȡ;�m}��,����-�� �
�����
�J�P   P   J�;�`@;�T`:x1��u���q�� ��'�����O������o�؞����n�� �PA)�_�v:�D;[�;/O�;P   P   s��;�G�;�`@;�
�M�����ż��S9�jg�+�����̓f�P-8�0���y��C�{����G;�q�;�[�;P   P   ��<t�<X6�<H�<���;;��^-�uP�s0��r9��3"˽�����Q��^$N���޼�� �28�;��<�9�<���<P   P   ���<��<鹱<ٿ<�M�;>�[�Y�$����������\$�`�>���>��#����^'���I"���S�H<�;���<z��<P   P   �9�<߽<�b�<��<L/�;�����M�q�ν�/�[���Ʀ������Q���񀾝�-���̽�J�����bэ;���<P   P   ��<Y�<xݦ<K`�<�?�;����a]�ד��[�(ӵ�6���''�u�&��������Y���CZ�����R<�;P   P   E8�;B~<���<r|<���;_�[���M�̙�%�m���ھ̔=�����^��򁎿�\<��@پ:�k���	�J���S�P   P   �� ��k<_Ij<$)i<���;4�M�$�IϽ2�[���ھ�0X��ɿÕ��/���ǿ��V��@پ��Y���̽�I"�P   P   ��޼~�,�S�<�@<t�
<M@����Ҝ�K!/�������=�X8ɿ_0C��z��AB���ǿ�\<�������-�['��P   P   V$N����E�:��<d� <�k�:Vw��~P�����Mǁ����h�����{��z��/�񁎿������P   P   �Q��K�
9�7�F;$��;'^?;���I�P�����$��'��ն'�F'����^0C�����^��s�&��Q���#�P   P   ����^�(��r���
���<;Ѝ9;w���%w�g*��Ͻ���?�����ն'�h��W8ɿ�ɿ����''�������>�P   P   ,"˽%�E��NIԻO�~��:����ٻt�zG�1̽��?��'�������=��0X�ɔ=�4��Ʀ�\�>�P   P   k9���F�<&���q���+�u'i� \���>2����庼zG��Ͻ���$�Lǁ�������ھ��ھ%ӵ�Y����\$�P   P   m0��ɪ)�E�����pf�[�����S��۵��m���t�g*�P�������J!/�/�[�"�m��[��/�����P   P   jP��P�)u�R�ջ��+��h���R���j���۵��>2�&�ٻ�%w��I�{P�Ҝ�FϽș�ғ�k�ν����P   P   L-�ށ�rB�Y��ދ���M�Z�K��R��X�S�[]�� �������Tw�����H�$���M��a]���M�P�$�P   P   ��[�=�֭�:9�B;��<;�.�:�M�5i��ኮ��+i���:��9;^?;�k�:M@�4�M�[�������!�[�P   P   ���;#
�;��
<L� <b��;��<;�����+��f���+���~�_�<;��;[� <s�
<���;���;�?�;t/�;�M�;P   P   %H�<��{<�h<�.@<E� <��B;�����ջ>��r��IԻ�
���F;��<�@<#)i<w|<Q`�<��<�<P   P   \6�<��<S�<��h<��
<+��:�B�Mu�Y���Q&��+�8�r�G9�BE�:D�<WIj<���<{ݦ<�b�<�<P   P   t�<g�<��<��{<�	�;��=�ށ��P�Ԫ)�F�1�E�i�(�^�����,��k<	B~<Y�<߽<��<P   P   ��,=�P)=�=r�=���<�_<�6&�ݬ
��km�y�������A��>�k����8��� <���<�f=�y=x�)=P   P   w�)=#`)=x�=�s=t�<]=�;|���:�p��ҽ�����.���.�m;� �нn�p
��Aj�;F��<JD	=�=P   P   �y=M�$==xr=i��<o�;��C������.r�,ϝ������h���p�U��k[��k����".;�G�<KD	=P   P   �f=wP="=�=�c�<��;�Q�2�ɽ&SJ��?������=K��������<���H��ǽ�E��".;I��<P   P   ���<-=Ĥ=M�=ٻ�<ᯤ;,"���ɽ�3\���Ͼ&;1�b&��|J������90�[�ξ2qZ��ǽf���Zj�;P   P   � <VE�<;��<;:�<\��<H�<�䳼�I���WJ�J�Ͼ:�H�ݫ�����<�w�����G�[�ξ�H�i[��g
��P   P   ���b</��<���<x��<�^<o'�O
q�����S���^1�Bұ���!�I�K��� �v����90��<��S���n�P   P   w���9�1�<U�<W�<���<���8b�
��3ҽ2_r��B��Hj������GL�H�K��<���������p���нP   P   3�k���b�թ�;�m�<څ�<Y��<
P�;��h���m����������ݗ������!� ��{J�����h��k;�P   P   �A���׼/Ǻ�<�I]<�~\<ж<kl�x�ټv,��$1/�.�����Gj��Aұ�۫��`&��;K�������.�P   P   ����	�������;�<�2&<�%<���;ݓ�}�
�����$1/�����B���^1�9�H�$;1�����*ϝ���.�P   P   s�����	��:#��Y�:B��;Zx�;�U�;Ę�;�s�:߁&�}�
�v,����1_r��S��I�Ͼ��Ͼ�?���.r����P   P   ukm���ؼ����I;�:���;���;��;硤;���;�s�:ޓ�w�ټ��m��3ҽ����WJ��3\�$SJ�����ҽP   P   Ԭ
��f�2պ�;V7�;t��;���;Ӌ;ޡ�;���;���;�l溡�h�a�
�M
q��I����ɽ/�ɽ|C��0�p�P   P   y6&�|�99��;�p<�<��;NZ�;���;��;�U�;�%<Ƕ<P�;���8g'��䳼'"��Q���l���P   P   �_<?�^<�4�<o"�<��]<�$'<߼�;V��;u��;/x�;�2&<�~\<T��<���<�^<R�<��;��;��;�=�;P   P   ���<���<���<oE�<��<��]<��<&7�;Q��;��;w<oI]<х�<Q�<v��<^��<޻�<�c�<r��<t�<P   P   u�=ɀ=?)�<ؒ�<kE�<g"�<�p<��;&:�:^X�:���;�<�m�<K�<���<::�<N�=�=|r=�s=P   P   �=��=+q=;)�<���<�4�<_�;,3պ�����:#�Z���_0Ǻ���;�1�<&��<6��<ä=#==z�=P   P   �P)={[$=��=ƀ=���<%�^<�997�f��ؼ��	���	��׼��b���9��b<NE�<+=wP=N�$=$`)=P   P   Ŕl=_ti=�_=O�I=J�#=A�<�'�;���8���{���_Z��L7��ӝ�D��;Rd�<q�$=�6J=�Z_=��i=P   P   ��i=<}i=��`=� L=H�"=vU�<�����4�>ḽӒ	���%�"�%�1	�����Na2��ॻ�d�<��#=l�L=�Ua=P   P   �Z_=�pd=_=�K=��!=B��<zpq��Ό���/�j�0Қ�|ѩ����p�i�Q���0��,�g��!�<a#=m�L=P   P   �6J=�X=ۃX=��I=��"=��<�c��Y���@����"j��	�_��Q����1���}?�,7���0���!�<��#=P   P   u�$=?�C=��K=�C=u�#=u2�<�Rq�����S�, ̾�(�Kn��%����m�	O(��˾V�Q�,7��#�g��d�<P   P   \d�<�"=��6=HJ6=ZT!=���<;��@�����@�	�˾�c<��I����̿xa̿�ə�;��˾�}?��0���ॻP   P   ~��;�5�<�Y=��!=��=%@�<x�;X�4�H��s樾��(�UW��d��-�KE��ə�	O(��1��P��Ha2�P   P   �ӝ��Uc<���<_=��=�X�<�^<i!���ȸ�?�j�Im��e�n��̿\��-�xa̿��m�Q���p�i�����P   P   C7��S�����<ߏ�<U�<���<�g�<�c׺T9�z�	��֚�+)��i���̿d�𿢦̿�%��_�����0	�P   P   [Z����o�&�<:�<[�<���<7�<3\<+�s�넽X&�����+)�e�n�VW���I��Kn�	�|ѩ�!�%�P   P   w���w��NX�:�,<�EW<�)]<V<�8*<�p�:|����L��X&��֚�Jm����(��c<��(�$j��1Қ���%�P   P   ��`��������:�;��<@�<�T<�
<>h�;O��|���넽{�	�A�j�t樾�˾- ̾���0�j�Ғ	�P   P   ��8��r��+�:5�;�m�;�}�;��;��;��;9h�;�p�:.�s�U9��ȸ�I����@��S��@���=ḽP   P   �t�̺�`<@f,<O�<��;�J;��H;��;�
<�8*<-\<�c׺j!��X�4�A������Z���Ό���4�P   P   �'�;{�_<�@�<n��<�W<;�<В�;ȄJ;h�;�T<V<1�<�g�<�^<|�;0���Rq��c��jpq����P   P   M�<ͽ�<}�<��<t��<*j^<2�<��;�}�;&�<�)]<���<���<�X�<$@�<���<{2�<��<L��<�U�<P   P   O�#=߀!=�=W=���<p��<��W<4�<hm�;d�<sEW<�Z�<U�<��=��=ZT!=w�#=��"=��!=M�"=P   P   R�I=�+C=�^6=��!=U=��<a��<f,<��;E:�;��,<&�<Ώ�<Y=��!=FJ6=�C=��I=�K=� L=P   P   �_=h{X=��K=�^6=}=r�<�@�<�`<�*�:����V�:��<���<{��<�Y=��6=��K=܃X=_=��`=P   P   `ti=�Pd=g{X=�+C=ڀ!=���<\�_<��̺ r�v������$�o��T��{Uc<�5�<�"==�C=�X=�pd==}i=P   P   $E�=;Џ=Tϊ=�4�=��Y=r=C�<�^C��O'�����ޚ��j����)&�	=>����<�=xZ=�i�=C�=?ݏ=P   P   ?ݏ=я=�4�=ܮ�=Z4]=��=�;�������ƻ�LC3��3�qR��������ֈ�;��=�^=��=�Z�=P   P   C�=��=Fʊ=���=/�]=v=7T]�B6���E�����خ���������������䂽-�<�g�=��^=��=P   P   �i�=�P�=*;�=�&�=e]=�=�&��v��DQ��p������/���/�����达�UP����q׻i�=�^=P   P   xZ='u=t�{=d�t=��Y=.�=�.[��Y��D�f��$� yC��G���ژ�C)��N&C������e�����<���=P   P   �=u.P=��`=��`=��O=��=<�;�����Q�龔�Y�����ܿ��ܿB���Y���辰UP��䂽���;P   P   ���<$=Y�;=��B=o;=P\=�A�<�����:(��~KC�E�����������C�O&C��达�����P   P   �<>��D�<�9=Q�=�x=��=}��<VuB��$������0��f%����ܿ����ܿE)������������P   P   �)&�R��;�0�<�e�<���<ܽ�<:��<ie�;I�&�[�{���/�������ܿ�����ܿ�ژ���/����rR�P   P   h����S"�C:<��<���<bg�<	֎<j�7<�$�ශ���2������/�h%��H������G����/������3�P   P   ݚ��IQ����V;�<�U<��<�A<��<3[N;�����o����2�{��2���KC���Y�yC���$خ�OC3�P   P   ����N����t�9�͙;��=;C�:E):��7;+ĕ;�I9����᷁�[�����?(��$�%龬p������ɻ�P   P   �O'��M$��U;��;�':�-�b�������lF:#ĕ;[N;�$�M�&��$������Q�K�f� DQ��E�����P   P   �^C��o�;�v9<l�<t�?;\�}�sk�u��ȅ����7;��<a�7<We�;buB��������Y���v��F6�����P   P   C�<���<�ɸ<Gۏ<�E<��':����}k������':�A< ֎<4��<y��<�A�<p<�;�.[��&�ET]� �;P   P   w=�=%=b��<V�<�]<د':��}�.�I�:��<Ug�<ҽ�<��=N\=��=/�=�=y=��=P   P   ��Y=]�O=��;=��=F�<V�<�E<��?;��':�=;�U<|��<���<�x=o;=��O=��Y=g]=3�]=^4]=P   P   �4�=��t=��`=�C=��=Y��<9ۏ<F�<��;c͙;�<��<�e�<I�=��B=��`=d�t=�&�=���=ޮ�=P   P   Uϊ=HC�=�{=��`=��;==�ɸ<tv9<�U;�n�9��V;�B:<�0�<�9=R�;=��`=r�{=*;�=Gʊ=�4�=P   P   ;Џ=Q�=GC�=��t=X�O=�=���<zo�;�M$�`���]Q��T"����;�D�<$=p.P='u=�P�=��=я=P   P   >�=ᝣ=8s�=�G�=��|=� 7=���<�:Y�ޮE��
�����ż��]�D��U�Y��<Z�7= J}=�b�=�}�=���=P   P   ���=��=���=襗=�O�=��5=T&<�*��Jݽ~�2��_���^��|2��_ܽ
8)�*+<(�6=C��=�ӗ=4��=P   P   �}�=c�=cf�=��= ��=�f1=�:cc��M>�혥��_�3���*�:H����=��K��/�}:c�2=���=�ӗ=P   P   �b�=�ؗ=�ȗ=�1�=\C�=j1=��a�t�ýs炾������D���w�_�w���D�g���9�����½�KH�d�2=D��=P   P   J}=�ω=���=��=�|=��5=�b':J�ýx�����n ����ǿMN⿤�ǿ9���z���4����½��}:-�6=P   P   a�7=�,h=�tt=mOt=��g=�7=Su'<pۖ�1�����dd���U �`�%���%�=] ��n��{��:����K��<+<P   P   i��<�I+=.�D=��H=��D=T�*=�T�<U�)���=�|W���Ŋ��< �Ĕ<�+
W���<�>] �;���k�����=�8)�P   P   �U���<�U=�s=`P=�
=�߼<#�V��+ܽ5����`D��Uǿk�%�B�V�-
W���%���ǿ��D�>H���_ܽP   P   Z�D���=;:�<���<췰<J�<<u�<p�8;shD���1�:x��v�m��m�%�ǔ<�e�%�TN�h�w��*��|2�P   P   ż��҉v�&J�;v�<�L�;k_�;ho<���;υv�v2��^��<���v��Uǿ�< ��U ���ǿ��w�3����^�P   P   ���"/Ӽܵ��a�8�={ϻ�L��ѻ�">�=v��ՍҼ�=��^�=x㾡`D��Ŋ�kd��u ����D��_��_�P   P   ���|Ӽ���4��<y��P�������bz�ԙ�ZA�׍Ҽx2����1�9����W��	���������������2�P   P   �E�x����<�gY��H=ۼN$����ۼ��ڙ�Nv��ۅv�yhD��+ܽ��=�6���x��z炾M>��JݽP   P   �:Y��)6;b��;�7�]�x�sۼӂ	���	�Īۼ�bz�#>�ౣ;.�8;=�V�a�)�yۖ�V�ý��ýmc���*�P   P   ���<��<f.�< z<��̻����X���ւ	�Y$������ ѻQo<2u�<�߼<�T�<<u'<a':V�a���:K&<P   P   � 7=.+=�d=?Y�<]��;��ƽ��ۼY=ۼ�P���L�%_�;J�<�
=Q�*=�7=��5= j1=�f1=��5=P   P   ��|= h=_�D=��=ζ�<F��;��̻��x�~Y���<y��{ϻ6L�;ط�<YP=��D=��g=�|=]C�=!��=�O�=P   P   �G�=?Ή=t�t=OYI=��=5Y�< z<v7�p�V4�Q�8�=�<���<�s=��H=iOt=��=�1�=��=饗=P   P   9s�=�ޗ=��=r�t=[�D=�d=V.�<��;]����O����I�; :�<�U=%�D=�tt=���=�ȗ=cf�=���=P   P   ᝣ=v��=�ޗ==Ή=h=)+=��<_)6;x��|Ӽ4/Ӽ��v�Ϥ=;��<�I+=�,h=~ω=�ؗ=b�=��=P   P   ۸�=v�=B#�=v�=,��=�*7=3;v<�gƼ?ʉ�3�ѽ�x�N?ѽ�W���ļf�x<��7=W̃=�r�=\�=�=P   P   �=��=�C�=��=�7�=@�@=M�;R�d�d �<�h������쑾�2h�:��$	c��m�;ЂA=�a�=��=�H�=P   P   ]�=v	�=��="��=*�=-#A=(�"�Z���_v�Iwܾ+r�6�/��T��%ܾ��u�Ag��U`���A==>�=��=P   P   �r�=BU�=�K�=�V�=�(�=i+A=1޻���������9.��f��)õ�޺���Q��>.��J�������Ի��A=�a�=P   P   Z̃=wl�=�p�=	W�=��=��@=���(e��U����\�<οZ&��d-�i&�1:οb�\�s�������6`�ՂA=P   P   ��7=;�b=��i=5�i=B�b=�7=��;΄���3��Hp\�ui��E�o-���3��U�E�h��c�\��J��Cg���m�;P   P   ��x<,�=:*=��*=9*=�l=`�w<��b��Ru�B�-��Ϳ��E������p������V�E�4:οA.���u�#	c�P   P   ��ļ�'p<)�<�,�<��<�ͽ<֝o<Vļ�8�)h۾~ی����M���AZ���p���3��m&��Q���%ܾ<��P   P   �W���=$��*z;��^;�n;"];�{x;�n#�����#g�Р�!����,�N�������r-���d-�溵��T��2h�P   P   Q?ѽc��/]c���y��d��ρ���`z�Gc�xH��н~!���/�#�������E���E�a&�3õ�?�/��쑾P   P   �x���8��ټ�1��w��FO*����h��?�ؼ��7���!��Ӡ��ی��Ϳ�i�!<ο�f��4r�����P   P   :�ѽ�9����������N���q���q���N���qW����7��н�#g�0h۾J�-�Sp\��\��9.�VwܾI�h�P   P   Eʉ��0�ټy����`�]��"施vp���&a�!��F�ؼ}H� ����8��Ru� 4��`���Ɣ���_v�m �P   P   �gƼ�X%��&c�0���ܤN�O��矡�㪡�wp����N��h��+Gc�o#�jļ��b�܄��;e������!Z��e�d�P   P   4;v<�Ro<U�|;{�x�v'�8Kq��˖�韡�&施��q�����`z�{x;��o<C�w<���;���s1޻�"��;P   P   �*7=$�=���<#lf;�Z����)�<Kq�	O��]����q�RO*�恟�w!];�ͽ<�l=�7=|�@=f+A=+#A=A�@=P   P   .��=!c=��*=	?�<);�Z��}'��N���`���N�����d��#n;��<2*=>�b=��=�(�=+�=�7�=P   P   v�=<��=�^j=_V+=?�<�kf;��x�I����������1��@�y���^;f,�<��*=/�i=W�=�V�="��=��=P   P   C#�=!r�=���=�^j=��*=���<͔|;�&c�ټ�����ټu]c��)z;�(�<:*=��i=�p�=�K�=��=�C�=P   P   v�=m�= r�=;��=c=�=�Ro<�X%��0��9���8�o��>$�l'p< �=1�b=tl�=@U�=v	�=��=P   P   ��=q�=��=Ή�=��t=LG=��;o3���½�}��p��Z�y7½#�2���;�U=�t=d�=�֥=�\�=P   P   �\�=d�=0��=���=.��=�n2=E:غ�3��Ռ4�=���t���}[���4�����Qo��·2=���=7��=���=P   P   �֥=QS�=�ۥ=|��=ӭ�=n�:=U$$�Y��l���m���H�K6c���H��?�� �����qw ��H;=���=8��=P   P   d�=���=���=�`�=Q��=��:=��f�(��>bվm`��E���p�g�9-��:`��վp� �c��H;=���=P   P   �t=H='�~=�A=�t=e�2=5�!�s����A⏿��
��}N��Hl��N�ۓ
��᏿���p�hw �ȷ2=P   P   �U=�9=L�9=��9=��9=�I=s̿�]����ԾԵ������!��DK�� S��=6�� ��᏿�վ���n��P   P   y�;F��<|��<�x�<Ǔ�<Թ<#L!;����#�����_��F
�)��x1��S0���M��>6��ޓ
�!:`�� ������P   P   �2�� ��L�ݹ�KK�sK�ѡԹ+�����1��S3�g�
��|��1�M���C!��T0��#S���N�?-���?��4�P   P   x7½�\�/sԼ-~����
�x_��Q�Ӽh���������^�G�	^�l�k���z1��IK��Il�g��H��[��P   P   �Z��x}��kH��h����������g�T�G�*'|��r��͵�B�a�^�5�M�,���!���}N��p�W6c� ﶾP   P   �p�*��������]��M�����ƽa����D��G9������V��͵�a�G��|���F
������
��E����H�~��P   P    ~�a���󠑽����߽ZA��A��r߽;��.J������r���l�
���_�ܵ��J⏿m`�n�E���P   P   ��½�}��~�����5��I��+�PK����<��I9��1'|�����S3�*����Ծ��Lbվl����4�P   P   o3�0i��;H�08��
�޽VB����
�QK�u߽�D��[�G�q����1�����o����5��m���3��P   P   z�;Sը�Q�Ӽ�g�6Z������!����+�
A��g�����g�e�Ӽt���K!;ο�x�!� �f��$$�\;غP   P   NG=�*�<�"���(���:���Xƽ���YB�	I�bA��ĕƽ�����_���Թ�ӹ<�I=_�2=��:=j�:=�n2=P   P   ��t=�N:=���<#�?��K
��:��:Z���޽=���߽X��������
�OK����<��9={�t=P��=ӭ�=/��=P   P   Љ�=:�="�:=�ھ<Q�?��(���g�78���������]���h�V~���LK��x�<��9=�A=�`�=|��=���=P   P   ��=f��=�&= �:=���<)&��e�Ӽ�;H��~����������lH�YsԼ��ݹ]��<A�9= �~=���=�ۥ=0��=P   P   q�=y�=f��=7�=�N:={*�<�ը�6i��}�e���/����x}��\�E!��(��<	�9=H=���=PS�=d�=P   P   �ޣ=bڠ=���=��=�fA=i��<����,<���e���3���F���3��:����#ɛ���<��@=ݚ�=�~�=���=P   P   ���=:Ǡ=t��=d�=�t=;
=��v�,�½�"S�d��0BѾm.Ѿ�馾-�R��A½�u�{�	=DJt=�-�=�e�=P   P   �~�=k��=�=�S�=쇂=Z�=�ɜ��y
�����A/���c�=����c�����b���"
��ʛ�d�=vf�=�-�=P   P   ���=�Ɂ=Ӂ=Ĵ�=ۂt=�=�:��V?*���"�}��2ֿK��Ę��ֿ�]}��y�*�L���g�=JJt=P   P   ��@=#IB=�K>=�mB=gA=�8
=�n����)����r������2n��L���4n����t������*��ʛ���	=P   P   ��<Î�<9��<�ɻ<��<�ŧ<�9s�/�	���>��)�5��k���������ˁ���5�t���y�"
�Śu�P   P   ɛ���y��Ի�o�L�һD�r��.��a��6٩�R�|�����H��P�������O���́������]}��b��A½P   P   ��������"��<�X�<���"�U��b:���Q�O��Hտ��m�������� �������4n��ֿ���/�R�P   P   �:��ᘽ�=���G���H���#��!떽�3���t�|����Ob�h�
��������R��������L��ɘ���c��馾P   P   ��3���ٽ�eսbs��	�	�{�	��6��G�Խ��ؽ��2�z�ϾLE��i�
�m��H���k��3n�R��D��u.ѾP   P   ��F�Z^ ��| ��'�'�0��9��0�����/ ����pE�{�Ͼ�Ob��Hտ���1�5�����2ֿͪc�:BѾP   P   ��3�` ��X��)�>�J�)�_�_y_���J���(�	�����2�����O�]�|��>�� s��2�}�K/�m��P   P   �e�!�ٽ�q �V)�PIT�0t����S%t�I4T���(��/ ���ؽ�t��Q�?٩���$�������#S�P   P   /<���Ř�4:սO�d�J��*t�������T%t���J����L�Խ�3��j:��a��9�	���)�d?*�
z
�9�½P   P   ����-C����&��[�0��r_�6��������cy_� �0��6��(떽b���.���9s�o���:�� ʜ�	�v�P   P   o��<�,q��"�ۭ�޹	��9��r_��*t�0t�/�_���9���	��#����"���r��ŧ<�8
=	�=U�=:
=P   P   �fA=r�<gE̻+�;���	�^�0�i�J�VIT�D�J�.�0��	��H��k�<���һ��<aA=ׂt=뇂= �t=P   P   ��=C=�i�<��.�;�ۭ�&��T�\)��)��'�qs���G��$�<��o��ɻ<�mB=´�=�S�=d�=P   P   ���=p�=Z?=�i�<�E̻�"�"���<:ս�q ��X��| � fս�=����"��Ի��<�K>=Ӂ=�=t��=P   P   bڠ={֖=p�=C=i�<�,q�4C��Ř�%�ٽ` �]^ ���ٽ�ᘽ����y����<IB=�Ɂ=i��=:Ǡ=P   P   �=]�=�et=@�?= "�<O��vL�Inٽ��*��H]���p��4]���*�`yٽ	M����1�<լ>=��s=�*�=P   P   �*�=�C�=��=�	o=�7=2��<S\�9��}�d�d'��1�ؾu�ؾ'����d�ё�ב�g<�<�66=�Gn=ܡ�=P   P   ��s=Q�s=t=�n=�P=ɒ�<�3��n�����A��I_���|��$_���� S��:�R뼆w�<PSO=�Gn=P   P   ެ>=��8=�9=�#?=��6=���<$��-�)��?羧�u��gϿJ<��6��LϿOxu��;{)��뼍w�<�66=P   P   ;1�<a:�<_Ϯ<p�<�b�<m��<���;P)�>#�۱����pif�s��sjf�n������*�;{)�R�|<�<P   P   ������ػ1=�`o<�-Ի񧷻�d����#�����Y/� ���#����¾�����[�/������:�ʑ�P   P   	M���3�7�U��bg��6U�)3�x�K��b�,����t�&N�&c���$��r���2:������q��Sxu�S��͑�P   P   Vyٽ����7Ƚ#߽y�޽��ǽU`���Lؽ�pc�7��ο�e�������s����¾�yjf��LϿ�����d�P   P   ��*�QG��w�6�'��0� �'�#+����S�)����(�]�����������$��&���x���6��$_�*��P   P   �4]�"�,��L=���\��q�-�q�s|\��<�r4,���[��'׾bB{�����e�*c��%���zif�P<�	�|�|�ؾP   P   ��p���C��pZ�����:����&���ゾ��Y���B�~o��'׾,�]���ο+N��Y/���hϿ!I_�9�ؾP   P   �H]�C�C���d�qx�������򷾐跾C|���K��]jd���B���[����<��t���䱝���u�J��k'��P   P   ��*���,�B_Z�$t��c~���iǾXо'YǾ�`���K����Y�u4,�X�)��pc�4���0��F#��?������d�P   P   Jnٽ�%�1+=�_���蒨�.iǾ��ؾ��ؾ(YǾE|���ゾ#�<�����Lؽ�b潘��GP)�9�)��n�C��P   P   vL�ǵ��zG�b�\�).����о��ؾZо�跾&��x|\�'+�]`����K�e���J��4�Z\�P   P   �N��t3��ǽ�'��q�����0iǾ�iǾ��#��5�q��'���ǽ93�U���Y��<{��<���<1��<P   P   ("�<�_ϻcT�~޽�l0��q�+.��뒨�f~�������:��
�q���0���޽7U��-Ի�b�<��6=�P=�7=P   P   B�?=�j�<k�8��`f�~޽�'�f�\�b���)t��vx�������\�?�'�3߽cg��o<�Z�<�#?=�n=�	o=P   P   �et=��9=�ְ<t�8�cT��ǽ~G�6+=�I_Z� �d��pZ��L=��w��7ȽQ�U�[1=�DϮ<x9=t=��=P   P   ]�=�(t=��9=�j�<`ϻ|3�̵���%���,�H�C���C�)�,�YG������3�<�ػD:�<��8=L�s=�C�=P   P   �vW=u�J=��"=s/�<���6�,����2�t\��0���㐾//���\�0Y�}}��A!.�:s�����<��!=�UJ=P   P   �UJ=ؚJ=�==�{=�}�<�iݻ'g�y����n�G��(ѾpѾ'���rn�C����g������<�_=�==P   P   ��!=)"=w"=�N=�Q =ya!<��$����.��L�J�?��W���?�6.�}��c
��%�v�<QO�<�_=P   P   ���<鰡<#6�<��<�<~�!<����i�`'ƾ��L��L��Qnݿyeݿ�7��1�L��ƾu�������<�<P   P   �r��cI(���V��	&�*J��KܻS$��-���پ�L������l�:���U���:�u���oP��_�پu���%�S��P   P   )!.�=N�GWo�o��M��,�0f�>t���ž�#��NK�9�t��˟��ҟ�&�t��l�pP���ƾb
���g�P   P   n}���˽.�r���k��5hʽ`u�����;v���'L��Y���Ut�Go��:�������(�t�y���4�L�~��?��P   P   )Y�ۥ��q5�\!G��G��5�!���N3m��������@:���������;����ҟ���:��7��8.��rn�P   P   �\�B�U���v�s�����7���]Rv�%U�T�Z�����>�sܿ�IU�����Jo���˟���U��eݿ��?�)��P   P   ,/��]F���K���ر�T����������������Ё�fy����Ͼ�kV�sܿ�@:��Ut�A�t�s�:�Znݿ�W�sѾP   P   �㐾�ˏ��p���3о�� )������Ͼ��KG��G����Ͼ�>� ����Y��TK������L��R�?�(ѾP   P   �0���Ǐ�H����,ᾎ��^��S�e��W�ྡྷK��LG��hy���������'L��#���L����L�L�L��P   P   s\��7���d���'ᾄ�	�(j�S##�X�N�	�X�����Ё�Y�Z�U3m�Av���ž��پk'ƾ�.����n�P   P   �2���U�\4��1%о��l���)�>�)�X�f���Ͼ����*U������Ft��-��i���|��P   P   ��I^�v�޿���뾋b��,#���)�U##��S�¿뾈���dRv�"!�ju��Bf�1S$�Ʈ���$�)g�P   P   0�,�*oʽ�5�񙋾����T1���b�l�+j�^�&)������;����5�@hʽ)�,�uKܻ\�!<ia!<�iݻP   P   ���VyL�j���F�!	��������!����	������[������G�x���M��J���<�Q =�}�<P   P   w/�<ٛ"�!�m�P����F�󙋾῱�6%о(��,��3о�ر�y���f!G�����'o� 
&���<�N=�{=P   P   ��"=���<�Q�#�m�j��5�ǋv�`4���d��N����p���K����v��q5�.�aWo���V�6�<yw"=�==P   P   t�J=q�"=���<�"�\yL�/oʽL^���U��7���Ǐ��ˏ�bF��M�U���˽XN��I(�Ѱ�<)"=՚J=P   P   ͼ=� �<��z<��$/�S$��N�nJ[�s�������'��i����1����[�������@1�Tj��u<Ҷ�<P   P   ض�<�f�<R��<�[<��Ļζ�׍��v�"�Q�|���d+ȾZ(Ⱦ���v�|���"��P����O�һ�V<֗�<P   P   /�u<�{<�x<�6[<�V�;��`��i�
��)Ň�Xwܾ-��&'���aܾ	Ǉ����j��g�B	�;�V<P   P   j�͆=�<�<.�h}ƻ�M`�6B�[��n�����s�����t���6�r����y��|����C���g���һP   P   *1�E	U���d��:T���/�����th�|M��¦���8�'m������c�a����p���8�����{���j�	��P   P   ���Tؽ���̪��j׽:	��?	��'����Q�8�\*ÿ"�%�>�Y���Y��&�Zÿ�8��y�����P��P   P   ����=.�� F�ŏO�<�E��-�i���"�@+��,����_�%�eIy�����xy��&��p����Ǉ���"�P   P   �[�jaw�熏��O��:���H��c�v�!�Z�e[{�0Y۾�r��!��wTY�َ�����Y�f���;�r�aܾp�|�P   P   �1��I����K��2�վ��޾��վ	��4�����i%��!W��������yTY�hIy�C�Y�g�x��������P   P   d����\���P�^����������,�徧����ǧ�ǾH9&������!��b�%�'�%����������&'�Z(ȾP   P   �'��aQξk����� ?3��";��3�����P���;P��Ǿ#W��r����c*ÿ.m���s�-�e+ȾP   P   ~����Iξd���+�'�J��]]��I]���J�^�*�]����;�ǧ�l%��6Y۾1�X�8���8�#��_wܾ��P   P   q��pE������+��]S��_q���|�C;q�7!S�^�*��P��������l[{�E+������¦�n��-Ň�R�|�P   P   jJ[�m���_2�S��˺J��eq�O��	��D;q���J����0���4��'�Z��"�-��M�b����v�"�P   P   �M���v�| ������?3�4l]�L�|�P����|��I]��3�����j�v�o��I	���th�6B��i�֍��P   P   O$��g�-�~Q��I�վ���3;�6l]��eq��_q��]]��";�����վ�H���-�D	������M`���`�̶�P   P   $/�_ ׽d�E�-&����޾����?3�κJ��]S�,�J�?3������޾:��E�E��j׽��/��}ƻ�V�;��ĻP   P   ���JS��ｶ:O�.&��K�վ���W���+��+����c��;�վ�O��ЏO�۪��:T�n.�t6[<�[<P   P   ��z<Q�7��c���f�E��Q��� ��e2澱��i��p���P��K��� !F���ｫ�d�=<���x<K��<P   P   � �<i�~<S�7��JS�c ׽k�-��v�q���uE���IξiQξ�\��Q���xaw��=.�eؽ^	U��=�c{<�f�<P   P   0oK<�U�;׾=�;�.����w����]��m��
Ż�d<׾�s�WN׾�껾&���r^�61��I����0��C�VC�;P   P   uC�;���;&S%��p��B ��|���7��XJ��m������ʾ��ʾ�'�������J����ݬ��>"�aEw����P   P   �C���6�� @�1�p�z`��X�.��U����k�v��{��Յ�����S��v���Tw��u��v���^1�Y�¼IEw�P   P   ��0�/�>��>��a/�r ���.��䅽~���|�t���Ծ)g �̐G��G�d ���Ծ��t�%����&���^1�0"�P   P   �I���a̽�ս�˽1L���\�����h��Y�w���S�Nc������|f��&&S�#/�Ôx�"����v��Ҭ��P   P   ,1�H�.��,>�R>�n.�\����������s�����i�&���t������C��j5j�#/��t��u����P   P   sr^����o���w��ލ��7���
]�%�I�׻u�%"Ծ<�R�����6���"����C��'&S���ԾOw��J�P   P   ���Џ��d ѾF��t��˦о�
�����mь�����������'���!��"�����f��d �t�������P   P   �껾k㾀��X��'H!������u��&��c5���M龝�F�:!��)��8���t�������G�S�꾀'��P   P   PN׾l��&���D�#�V��V��D�'G&�i��]־�ɾ�o����F���������&��Rc��ѐG�������ʾP   P   �s�'��1<���h��v��:ڋ��W��Xsh�a�;�Q9�z��ɾ�M龢��A�R���i��S�-g �؅��ʾP   P   ^<׾����D�=~�gM���M���:��@���}���C�R9�]־e5�����+"Ծ�����Ծ�{�����P   P   Ż��[�H'<�l~�/֠����(�ſgZ�������}�c�;�j��)��qь�޻u���s�b�w���t�m�v��m��P   P   �m��Q7��&���h�XQ�����F�пJ�пhZ��A��[sh�)G&�y�����+�I���#h���������XJ�P   P   ��]��M�������D��{��U_��c�ſH�п*�ſ�:���W���D����
��]�������䅽�U���7�P   P   u��|ł�w�о2����V��틿V_���������M��=ڋ��V����Ҧо;���c��]����.�[�.��|��P   P   ���{�-��}�����G!���V��{��[Q��3֠�kM���v��*�V�,H!�|��䍓�v.�<L��r ��`���B �P   P   :�.�oZ˽�=�ؙ����3����D���h�s~�E~��h���D�^��O��~��\>�%�˽�a/�T�p��p�P   P   ܾ=���<�$ս�=��}��z�о�����&�M'<��D�1<��&����m Ѿw����,>�.�ս�>�� @�4X%�P   P   �U�;K�2���<�qZ˽~�-�ł��M��W7��[����,��l�k�ُ�����R�.��a̽C�>���6�y��;P   P   	�뻠�r������ y
��V�뗾Ⱦj���Á
�#x�I�
�O���)OȾ�B���V�R'�('���%�N%v�P   P   ;%v��Et���ü�)0��|�����I6�
O�d禾.~ɾ�2޾�=޾��ɾ��������6��\���И��H2�zkƼP   P   �%��_�\!��_0�L�\�"���g��2q*��4v��O��\5Ⱦ��վ`EȾ�t���v��+��$彵���v_��H2�P   P   '��D2���觽9S��-�������ڷ���x�N�L}���ؾ3� �p� �$�ؾ[���r@O�����x������И�P   P   I'�����v����݈
�V��XN���:D�x�������)��<�})������
��{�D����w$彃\��P   P   ��V�"Ww��r��EX����v�6�U��5�,�)�Q"N�7���(2��J�s�}�4�}��EJ�Cl��
��n@O��+���6�P   P   �B������˾" Ӿ�ʾ��������;�~��>u�#��;����I�Ty��N���ږ���EJ�����Z����v����P   P   OȾ�����E�JV��?�1�����Z|Ǿ]@��5���/ؾ"�(��'}��|��O���6�}�~)�#�ؾ�t�����P   P   D����#�N'=���V��m`���V���<�å����R�Ⱦ�/Ǿ�H ��t;��'}�Vy��w�}��<�p� �\EȾ��ɾP   P   D�
�%K6�.i�����0���|���9w��j�h�<�5���	��ݾU�Ծ�H �$�(���I��J�)�4� ���վ�=޾P   P   x��F�������ſ��пφſ��������VE�@���ݾ�/Ǿ2ؾ�;��+2�����ؾZ5Ⱦ�2޾P   P   ��
�� F�j<��0���������ˊ�����Պ��VE���	�U�Ⱦ8���&�;���|���N}���O��*~ɾP   P   c����56�������'>��^R��� �*�,����������>�5����`@���>u�V"N�?D�{�N��4v�`禾P   P   Ⱦ��@i���r���Z�y�,��,�*�͊����n�h�ƥ�^|ǾB�~�1�)�����1q*�O�P   P   뗾N5���=�h���}�ſ�)�r!�{�,��� ���Ԇſ<w����<����������5�`N㽹ڷ�f��F6�P   P   �V������!�9�V������ѿ�)��Z�aR�����п������V�6�Ċ��>�U�a�����$������P   P   y
�7�v���ʾ�@�Dw`������ſw��->����鿆�ſ6����m`��?�"�ʾ��v��
�5���S�\��|��P   P   ����N�+/����Ҿ�@�;�V�j��������7���󨿌�����V�QV�+ ӾKX�����DS���_0��)0�P   P   ���K����+/����ʾ�!��=�Fi����o<�����%.i�W'=��E��˾�r���v��觽j!���üP   P   ��r�6?��K���N�9�v�����S5�����56�� F��F�-K6��#��������/Ww����P2���_�Ft�P   P   	�����*;}�0���8:����8�þ����D���/��H7���/�п�T����&ľBn���:�����z��P   P   u��b��e6������۽[�$��/k�������Ⱦ@^�S� �4� ����q�Ⱦ�����l�D}%�ܽ�ȍ�=�7�P   P   ��Nv���}�޳��zD��!۽�:��I�㮅��T���{��.~˾I�����������J���ܽ�����ȍ�P   P   }��h���Q뽻�㽢$۽�۽z�� ^�M�E�])���p���Ἶ�＾�����q��g_F��G�Hw�
�ܽ��ܽP   P   
�:��L�naR�v�K��=:�|�$��=/�'0��]m��d���"ɾ	�پ�Eɾ-���1)n�u#1��G� �<}%�P   P   :n���Wj���I��	E���㋾\�j�KPI�E�cm�����eپF� �� �ޱپM���/)n�b_F���J��l�P   P   |&ľ����������k�Zaþ���-������]���)پ=|
����V�
�ޱپ,����q��� ������P   P   G���W�'�:��
K�`�J���:����/�����Ǿ����س��q}Ⱦ�� �!������ ��Eɾ����ڌ��h�ȾP   P   ɿ�K��O{�c$����������z�qJ�(�CP�z{��b���M�ؾ�� �>|
�G� �	�پ�＾C���}��P   P   ��/�9�p�4<���¿��ؿ��ؿ�����ǝ�,�o�./�a����^ʾc���r}Ⱦ)پ�eپ�"ɾ�Ἶ)~˾/� �P   P   �H7�B���ٷ��-����/-���3��=��7���|6�b���{{��ڳ��_�������d���p���{��N� �P   P   �/�����-���Ə	��[5���S���S�D�4��'	����8��0/�EP뾅�������gm��]m�])���T��9^�P   P   ?����p�ҷ�Z�	�"�C���z�؈�5?z��4C��'	��=��/�o�*���Ǿ-��E�'0�M�E�அ���ȾP   P   ������J��.��9/�ch5��z������8?z�G�4�8���ǝ�	qJ�5������PPI�@/� ^��I�����P   P   4�þ�'�O,{�`¿���S��������؈���S���������z����_aþc�j��}���:��/k�P   P   ������/�:�s��p�ؿ�X���S��z���z���S�5-���ؿ������:�k��㋾��$��۽!۽Y�$�P   P   �8:�#D�������J��'��q�ؿ�gh5�)�C��[5������ؿ��h�J����E���=:��$۽D���۽P   P   0��nK��"��� ���J�t��c¿?/�_�	�ˏ	��-�¿j$���
K����I����K����峌�����P   P   ,;}���꽒�Q��"�� ��1�:�T,{��.��ҷ�4���ٷ�;<���O{�/�:����`j��yaR��Q���}��e6�P   P   
���u����nK�$D������'���J���p�����G���D�p�K�W��������L�v���Nv�b�P   P   �z���>�>�����`d�p���5����>�MX�
�a�eaX���>�'���ા��d�������� �?�P   P   �?�`�>��3w�e���L�	�B�J�ŧ���ҽ��|��
��1�;�Q�
� ��<�����8�K���
�Vŷ���x�P   P   ����r䟽^���������ٽ[�	�-�4�@7l�J��W��o̾1�Ծ�8̾WO���l���m�O�5�W�
�h:۽Qŷ�P   P   ������K���8�	���	�F	�^�)�gVN�{�|����������̢��ꔾta}�=O���*���T�
���
�P   P   ��d�Nx���,�w��d�̿J�7C4�_^)���0���K��(t�����'=��'�	�t���L���1���*�I�5�/�K�P   P   �ાc�¾Ġо�yо�a¾\=��x[���k���M��K���d����/�����Y����e���L��<O�zm����P   P   ���L�����B&�v���i�%��>���y��Y�{��is�څ��0���Y��t���Y���t�la}��l���<��P   P   '���D��|h���}�u�}�Fh�E,D��ŏ�1��q������唔��.���Y�����%��ꔾPO�����P   P   ��>�Q�~�BV��������Ŀ�W���럿$�}��>�y

�K�ʾ�ԡ�����攔��0��.�%=���̢��8̾K�
�P   P   [aX������Ͽ�������6�Y3Ͽ@w��t]W�go��zӾ�ԡ����څ������������*�Ծ;�P   P   �a�:ɨ�PA��c,���X�*lk�STX��x+�nJ������`�go�L�ʾr����is���d��(t�����i̾�1�P   P   MX��è��r�_�G��o���/�����q��q;G�A�����u]W�z

�1��]�{��K���K�w�|�R���
�P   P   ��>�����9����G����<}��B���S)��Y���s;G�qJ��Bw���>�ɏ��y����M���0�eVN�G���|�P   P   ����f~�a�Ͽ�,�k}������V���+��U)��s���x+�^3Ͽ)�}�	��>���k�b^)�^�)�<7l��ҽ�P   P   �5��D�ZC�����J�X��[��g����V��F������ZTX�
6��럿J,D�,��|[��;C4�H	�,�4�§��P   P   p��o��%Sh��������o�k��[�����C}���/��4lk����W��Nh��i�b=��ӿJ���	�[�	�?�J�P   P   ^d��m¾�����}�S�Ŀ���N�X�o}������o����X������Ŀ~�}�|���a¾�d�>�	���ٽL�	�P   P   ��ow�VYо~1&���}���������,���G�i�G�l,���������}��B&��yо7�w������h���P   P   ?����O�`�~�WYо���(Sh�^C��g�Ͽ�9���r�\A����ϿIV���|h���͠о��S��g����3w�P   P   ��>��F���O�ow��m¾q���D��f~�����è�Bɨ����]�~���D�S��l�¾[x����{䟽i�>�P   P   Q\5�>�f��ܿ�wu"������¾�		�'�4��	_�K|~��%���~�(1_��5��B	�*Nþ4j���#�c����g�P   P   �g�y$g�,���6�ӽ�W���g�6����fؾ�P����"+�-+���q}���ؾ~2��'�h�8)��?ս�T��P   P   [���3p���$��^	Խ���jb��pM�k������Ȩž��ܾ����ܾ��ž���m+���sN��[��7���?սP   P   �#�:w&��D&�O�"�SJ�>J�NM'�� <��#\�� �������B���V��Rޒ�r����]��==��r(��[�2)�P   P   .j������␾�Ì�e�E�g��M���;��8�XC�/�V�NWi��q���i�5�W�XD���9��==��sN��h�P   P   !Nþ��޾U�/(�n޾ޔ¾NZ���N��*�[���B�<>�ٿE�]N�}JN�@cF��A?� XD��]�h+��v2��P   P   �B	���$��R9���@�D9�V�$�"����׾�r�����KV�=_E�%D�p�E�7�D�>cF�0�W�m��������ؾP   P   y5���f�����d閿,Ζ��@��A�e�
P4����ľ"ۑ��4h�_M�fE�o�E�zJN���i�Mޒ���žk}�P   P   1_�ї�,ÿ���:������¿�8��� ^�?�_`۾�N��Өo�_M�$D�[N��q��V����ܾ��P   P   ��~�󓹿�t���*�t%F�Q�E��*����	����I}��9*��㾤N���4h�=_E�׿E�IWi��B�����,+�P   P   �%��	�ο]���Ei�`���R��A��Gih��,���Ϳ�y���9*�``۾#ۑ�LV�<>�+�V������ܾ�"+�P   P   B|~�3�οI�*�6���W+���_���#�����_��(�)���Ϳ�I}�?��ľ �����B�XC�� ��¨ž��P   P   �	_�у�������J1���w�ۆ%�t:�x��_���,����� ^�����r��-�[��8��#\�����P�P   P   "�4�>���_n�}Qi�{B��ͅ�q�5��5�v:����Lih�����8��P4���׾�N����;�� <�h����fؾP   P   �		�m�f�tÿg�*�?������3�%�r�5�ކ%�$��F���*� �¿G�e�&��SZ���M�PM'��pM�3���P   P   ��¾��$�Lu�����SF�B�������Ѕ��w��_���R��Z�E��濙@��[�$��¾M�g�BJ�kb���g�P   P   ��G<޾-9�薿`���SF�B���B��S1��a+��`��~%F�E���2Ζ�K9�w޾j�XJ�����W�P   P   wu"����5�J�@�薿��k�*��Qi����>����Ei���*����k閿��@�9(��Ì�W�"�f	Խ9�ӽP   P   �ܿ���%�خ��5�-9�Nu��xÿcn���R�*�f���t�,ÿ ����R9� U��␾�D&��$��0���P   P   A�f��׹���%����I<޾��$�r�f�C���؃��<�ο�ο�����ї���f���$�ǝ޾���Cw&�<p���$g�P   P   �a�g#��"�ֽm=0�󋾴gҾm�$�F���v�	����������� w�b�F�\J���ҾtT����0��l׽����P   P   ����=Q���}���%齣�*���x�I���=�龍����+���:���:�K,������pp��s�y���+�`�iD��P   P   �l׽K�ѽ��ֽ�.齍���)��4[��W��Ġ����Ѿɢ�q����PҾG��э��3\�p�*����`�P   P   ��0�!%5���4�{H0���*��)�|�1�#F���d��3��"��ʠ��ڵ���_������*�e��DG��3�m�*���+�P   P   nT��x��5N��P×��؋��zx�m�Z�g�E�f=�n�@�܋K�2V��)[���V��EL���A�x�>��DG��3\�i�y�P   P   ��Ҿk����Z��X�Ҿ�����匾Rd��p@���-�C�'��''�b`'�k(��
/���A�#�e��Ѝ�hp��P   P   UJ��S4�.TK���S�^
K���3������辡ޯ�󘃾N�J�a^'���p3�?5�k(��EL�{���?����P   P   X�F����/���H���Dv��rd��n�~�)�E����о�I���NU��o&����o3�_`'���V��_��GҾ���P   P   � w�_ժ�J�߿*���������޿m��o�u��+��B�4���׶Y��o&����''��)[�Ե�����C,�P   P   ����O�ӿ|6���M��,s�*�r��KM�m��$�ҿ����Xx9����4����NU�a^'�@�'�,V�Š��q򾟏:�P   P   �������^>��R���V���&��%���}���3c=�ã��Ǔ�Xx9��B辒I��O�J���-�׋K�"����龥�:�P   P   ���{���M��Z��^����v���j�{����L�ţ쿍����+�
�о�����p@�k�@��3����Ѿ��+�P   P   ��v���ӿ*]>��_��Z�>���O��=���}���5c=�'�ҿs�u����ޯ�Ud�f=���d��������P   P   �F������2��]�����M%>�� b�	 b��=��j�����q��q��-�E���辋匾i�E�#F��W��7��P   P   i�2���߿��M�����m��m�O�� b���O�z��+����KM���޿t�~��������r�Z�}�1��4[�F���P   P   �gҾ6#4�����h�us����n��P%>�>����&��6�r����wd����3�%Ҿ�zx���)���)���x�P   P   �;��5K�ٞ��{�us������`�d���V���,s����Kv��f
K��X�؋���*�����*�P   P   m=0�𻗾��+�S�ڞ��j���M��]���_���Z���R����M�1�P�����S�_�V×��H0��.齡%�P   P   #�ֵֽ4��"�����5K�������߿�2�2]>��M��^>��6�V�߿6���7TK��<N����4���ֽ�}��P   P   h#���Mѽ׵4�񻗾=��9#4�8��������ӿ������Z�ӿhժ� ���S4�v����)%5�T�ѽAQ��P   P   �N��x˶�`���|<�������׾(O�zM��{����������"��대��M�J~��ؾ�搾W=�����.��P   P   �.��b�{ͽ����2�(J~����ė�l��l1��t@��}@�:"1�S�����x����@�3��W��*νP   P   ��������.��q��}	�~-��
]��K��WI��aHԾ}�쾕�����ώԾ����|���E�]�d.�/���W�P   P   P=�~�C���C��z<��2�^Y-��2���D��~b�m���0�� C��pW���P�����qc��F��3� d.�:�3�P   P   �搾U������zٝ�Kk����}�ݑ\�O�D�vU9�u�9��A�-BI�d�L�ݠI���A���:��:��F�>�]���P   P   �ؾ���&Y��?������?׾v����̍���a�GI9��U!�������>���s�~i"���:�qc�w���x��P   P   C~�3a:���R�]�[�ŒR�V�9�������u�����>@�dc�0O��Ʀ�Sc���s���A������������P   P   �M�<��h!��sf���A������������L�x��OӾW/��>H�
��Ħ�;��֠I��P��ƎԾL��P   P   匀�������t��)���Q���쿮ⲿ���0��h�i.���PK�
�-O�����]�L�jW����2"1�P   P   �"��|��%��a��څ���� L`�G$��l߿
J��\N?�cM��i.��?H�dc����&BI��B�������}@�P   P   �����l���'O��ڠ��G��ދ��N���m)��NN���������]N?��h�X/���>@��U!��A�,��u�쾍t@�P   P   ����h����`������j�a�.�Ĺ.������f{_�����J���0�QӾ��HI9�r�9�i���ZHԾf1�P   P   �{��B��)O�_������[Q�>�c�aQ��o����QN��l߿��z��u����a�uU9��~b�RI��g��P   P   �yM�����|%�����~�nQ���v�ކv�cQ���p)��G$��ⲿ��L�����̍�Q�D���D��K�����P   P   %O��'����E!a�ف��y/�J�c���v�B�c�ȹ.�V���L`���쿶������z����\��2��
]����P   P   ��׾(9:�������'
��F��{/�nQ�[Q�g�.��������Q�����[�9��?׾��}�aY-�~-�%J~�P   P   �������Y�R��x�����)
��݁���~�����j��G���څ�0���A��̒R�����Pk���2�	���2�P   P   |<��ݝ�MF��\��x�����K!a���h��������ڠ��a�{��zf��f�[��?��ٝ��z<�t����P   P   `�����C��ڢ�NF�Z�R������%�)O���`��'O�%����p!����R�+Y�������C��.��{ͽP   P   y˶��M����C��ݝ����+9:��'������J���h���l��������<��<a:����\����C�����e�P   P   �,�N���&&���R�d����Ӿ==�TH���z�Ө������⯐�v�z�B:H�$c�4ԾMa���HS�qr&�V��P   P   V����G��=q�PW?�!�|�����:x�$��P�+�O;��&;���+�����������}���?����h��P   P   or&�<�)�8&�Ho�s`���/���U�Lȇ�E9���w˾����������˾���C,��3�V�`�0�N ����P   P   �HS�li`��?`���R�\/?�X�/�M�,��9�+�S��t��v���h���{��_�����u���T�Z�:�	�-�]�0���?�P   P   Ha���<��F$��1���g�g|��[U��29��@+���)��0�xU7��:��7�5�0���*��u,�W�:�,�V���}�P   P   +Ծ?�����%}�[���IӾ���`B��S!S��z)��D��u�A/������8��O���*���T�>,�����P   P   c��R6���N�� X��N�W�5����$|�>\��s�s��//�Q�ֽ$Rǽ�!׽6�0�0���u�������P   P   9:H�?'��+�������ы��
M��n���6>G���8?ʾȋ��=6�����$�ƽ"Rǽ�����7�Y�����˾���P   P   k�z�	���'O近V����J�翖Ү�4ly�>�*�;8�KP���	9�����ֽ;/���:��{�������+�P   P   ܯ�� �ۿF!�)![��2��5��mkZ�W ��_ڿdԏ���9���LP��=6�P��u�qU7��h�����&;�P   P   �������e�I��2��.���=���3q��炛��H��5��/����9�<8�ɋ���//��D��0��v�����G;�P   P   ͨ������Z�A���+���)���)�տ�Y��L�Y��5��eԏ�@�*�:?ʾu�s��z)���)��t��w˾J�+�P   P   ��z�h�ۿY�I�����U���K��]�}}K���Z���H��_ڿ7ly���@\��U!S��@+�&�S�@9����P   P   OH�×��!��E��wA���K�1�p��op�}K�׿�낛�W ��Ү�9>G�(|�bB���29��9�Iȇ�4x�P   P   :=�9��DT��E[��)��-2*�&*^�3�p��]���)�9q��tkZ�Q��q��� ������[U�M�,���U�����P   P   ��Ӿ�56������n�f����.2*���K���K���)�F���;����M��\�5��IӾ�g|�Z�/���/��|�P   P   b��h����N��ˮ�/H� f���)��zA��U��+�8����2���؋���N�c��j_/?�s`�NW?�P   P   ��R����*���X��ˮ��n��E[�F�����J���2��5![��V������ X�*}�6�����R�Io�<q�P   P   �&&�� `�S��+����N�����IT�!�b�I��Z�o�I�N!�3O�2�����N���L$���?`�8&�G��P   P   N��<�)�� `����h���56�<��ȗ��p�ۿ���"����ۿ���E'���R6�H����<��qi`�>�)���P   P   ��������K��t���뙾��ʾ�@
���7��Ie�"����������[e�k�7�h\
�x�ʾP��փ�Zc�����P   P   ���^���I~���d�D�_�J5~�ӡ��rӾKB�,=��N+�`T+��M��[�m�Ӿw����~���_�e�On~�P   P   Zc��v��VS��V�d��NF�)/;��JL���w�*홾�X����ξua׾�ϾՋ���3��_�x�X�L���;�Q�F�e�P   P   փ��ސ�vА�����m_�N;��'��k(�@�;���X���t������&Pu�P�Y��<��C)���'���;���_�P   P   L��%
��0�!خ�}���9�}�M�K��(����}���J����!�*!��r�c]�o���C)�R�L���~�P   P   p�ʾ(D���s�7��}ʾAE����v�U;���F��)�۽�ҽNӽ5�ܽ?���a]��<�V�x�q��P   P   c\
�w�)�TRA�� J�o
A��[)�u�	��yҾ����W�����ڽ����;���$���2�ܽ�r�H�Y��3��d�ӾP   P   d�7���n�kX��p���v��� ���m���6����'��M&s�����1ѽW��9���Hӽ$!�Pu�͋���[�P   P   �[e�é���>ѿ6�������Y��.�п�잿d�fE�ƃ;"ま5z ��1ѽ�����ҽ��!�����Ͼ�M�P   P   ����ƿ���p�>��^`��`�.%>�!+��ſ2H��J/*�~�վ"ま�����ڽ$�۽D����ma׾ZT+�P   P   ~����l޿O�0�5X��H�������>N���Ą�o�/��ݿ�ʉ�K/*�ǃ;N&s���C������t���ξ�N+�P   P   ��`l޿�y>��>������'4�j����p���[=��ݿ2H��hE�'����W���}���X��X��&=�P   P   �Ie�Dƿ֐0��F�����U.�r?�
.����p��q�/��ſ
d������W;����<�;�%홾GB�P   P   ��7�����?��kj��&����h.�|�P���P�
.����Ą�$+��잿��6��yҾ��v��(��k(���w��rӾP   P   �@
���n��Iѿ��>�����e��D?�~�P�u?�m�CN��4%>�3�п#�m�x�	�DE��O�K��'��JL�ӡ�P   P   }�ʾ��)�K^�����a�`��,���e��h.��U.�+4�����`��Y��� ���[)��ʾ<�}�M;�&/;�E5~�P   P   뙾���UA�ն�� ��b�`����,���������P����^`�Ʀ�v��u
A�=������m_��NF�@�_�P   P   s����设��%J�ն�������>�oj���F���>��;X��y�>�A���v���� J��s�$خ����T�d�~�d�P   P   �K��cĐ��綾���UA�M^���IѿC��ܐ0��y>�W�0�����>ѿqX��[RA��3�wА�VS���I~�P   P   ���{��dĐ��设���)� �n�����Jƿil޿m޿�ƿʩ����n�~�)�0D�)
���ސ�v��]��P   P   �k�����.���"/����¾ġ��'���gE�Rgb�@Wm��lb��qE����������¾\I���ļ�)����P   P   ��
���Κ��ה�k�Gd��������������r�b��群!������<懾�딾����7��P   P   *��-������7����Y��.�]�u�I�g]��Ä��Y��]4������H����������|]�cFJ��2^��j������P   P   �ļ���־"�־͸��V˔�n�]�(e+����� �7�6�x O���^�S�^�MnO�j7��� ��%�Y�+��2^��딾P   P   YI���";xپ;���&���=cI��4��#�����?������7�*^�����^e�>����%�_FJ�:懾P   P   ��¾9��y� ��� ���龈'¾T╾�\��S�kｈ�½�߮��:�������C�ĽYe�}� �|]�|���P   P   ��������.��6��.��g�����Q��	����a5�����X!��Sr���w� Z������d7������!��P   P   ���\-O���y��~��tc���x�NjN����h��>���sM����P榽Kcv��w�����%^�EnO�������P   P   �qE������x��T�ϿL+ܿ�DϿ�宿`��<TD�f��ٰ�8�\����P榽Qr���:���7�J�^��H��]��P   P   �lb�{p���n�|��/�E�.�h��p�m���ka��	��2��9�\����W!���߮�����^����l�P   P   8Wm��u���_��L�����g������/PK�q���h��h�k��	��ٰ� tM�������½7���q O�V4��~�P   P   Kgb��u��$T�`q��8���������歭���o�ڂ��h��la�g�	>���a5�k����1�6��Y�����P   P   �gE��p��ue�U*q�^ܿ��� ����Ǚ ��)����o�s��o���>TD�j��
����S��#��� ��Ä����P   P   #������~��;L�LV���� �HU�8�ș �譭�3PK��p�`�����S���\��4����a]�~���P   P   �����(O�b������g�����]'�IU�����������l��宿RjN�����U╾<cI�%e+�p�I�Cd��P   P   ��¾����y��ϿxH/��������� ��� �!����g��J�.��DϿ�x��g��'¾&���j�]�(�]�h�P   P   /��+����.�&�����ܿyH/�i��PV��cܿ��8������/�S+ܿxc���.��龾��S˔��Y��ה�P   P   +���Y;S� ���6�'���!�Ͽ����;L�^*q�jq��L�|�\�Ͽ�~���6��� �;ʸ��3���ʚ��P   P   ��`�־��ؾT� ���.��y�e����~�ye�*T�`��n鿿x����y��.�|� �yپ �־������P   P   �����b�־[;.�龐���(O�����p���u���u���p������d-O����?���";��־*���
�P   P   �B�������Q��o�i"۾��¾�)ؾK��.!���7��(@�ϧ7��2!�&��A:ؾþ7'۾hl���P����P   P   ���������`�'q"�t�ܾ����^Џ�d����\���m߾C����{߾�r�����⏾����Zsܾ�Z"�h�`�P   P   ��P���d�wQ��x"��%�@��ɚX�upG��J^��T��̫������ܹ���n��&�^�>�G���X��8��y�߾�Z"�P   P   jl�i�-�u .�����ܾf7����C�Ğ�����/�>)�{�6���6��x)������� ���C��8��[sܾP   P   8'۾x
�ŧ�Q�t۾jڟ�m=X�m[��iؽ-���x�ǽ7�ս��۽��ս��Ƚ�½��ٽ� ���X�����P   P   þ�/���iy�]��ݡ¾�e����F���G��ꚽd،�ú��3��[����X����½��9�G��᏾P   P   ;:ؾ�����I�$������k׾�Ԟ�M�\���nƽ�+����]���L�:c_�Y�����Ƚ����^����P   P   !���,���N��>c�c�
CN�_�+�=�P2���Y���'�1xӽ������K���L�/����ս�x)��n���r��P   P   |2!��Z[�FD���f���<��x$���֊��dZ�YI ���ݾcz���5���ٽ������]�������۽��6�׹���{߾P   P   ɧ7�}���n�����/�������L�m����e��ˋ6�%b������5�2xӽ�+��a،�0�սt�6�������P   P   �(@�ّ���Կ@����4�kC�c�4�EB��ӿ���,�>�&b�dz���'�nƽ
ꚽr�ǽ>)�ǫ��;�P   P   ��7��ّ��ῦ�'�Yf�#��m ��-te��'���࿱��̋6���ݾ�Y����F��(����/��T���m߾P   P   .!�k��֡Կ/�'��z����Z���w���l�y��'��ӿ�e��[I �R2��O�\����iؽ����J^��\��P   P   H��J^[��{�����j=f�b���������x���/te�GB�p����dZ�>��Ԟ���F�k[����opG�`���P   P   �)ؾ�,��P��
⿨ 5�aR��������\���p ��f�4�L��֊�b�+�	k׾�e��i=X���C�X�ZЏ�P   P   ��¾��%�N�0��� ���C�bR��d�����#��kC�����|$��CN� ��ܡ¾gڟ�a7��@������P   P   e"۾Q!� ���oc�Ɓ�� �� 5�n=f��z�_f���4�6����<��c����\��p۾��ܾ�%�o�ܾP   P   �o�) ��}�v�$��oc�2���

⿲��3�'���'�E������f���>c�K�$�iy�O����x"�$q"�P   P   �Q�c�-����}���'�N��P���{��ܡԿ���Կ�n��JD����N������ç�q .�rQ���`�P   P   ����1�d�d�-�* �T!����,�O^[�o���ّ�#ّ�����Z[��,�
���/�w
�f�-���d�����P   P   ����V���|q�W��O�Ѿ:\��3@־�^���m����m��_���B־M^��`�Ѿx���q������P   P   ������PԿ�5��ˡ)�މ;�x��ȑ��\@�������������[H��x���"q���g;|)����U/ԿP   P   ���տ���s@��ތ3���Ӿ�%��|�>�� ;�Z$S��ql�3�v�I�l��?S��=;��>����tXӾO3����P   P   �q��ˑ��ّ�Nq���)�ҞӾ�\w�K&�##������}�e��r����}�������>��1w�tXӾ|)�P   P   y��x�<�w�L��<�+���;6	�����\˽mZ���ҭ�ʹ����ý��cn��C(��<�˽�>�����g;P   P   `�Ѿ;��c��c��6�^nѾ�/����=�3�ʻ�����Q���O���\؇��Q���5��A(�������>�!q��P   P   J^���*���#���L�����9Ͼ���@�9�^'���������vTh�\�_�6�i��Q��_n��~}��{=;�t���P   P   �B־AD�7W'�o�7���7��'�s�
�2AվJ���xQ��0��躽����_�Z�_�Y؇������?S�VH��P   P   �_����)��[T���t��}���zt���S�@�(������̯��jj���O�������uTh�L�����ý�r�A�l���P   P   �m�>H��L���硿�B�����;���҃��EG����ְ���t����躽���P���ȴ��e�,�v����P   P   ���W[�Qo���ɿ�y�� �5�jȿ_̘�u5Z����ְ���jj��0���������ҭ��}�zql����P   P   �m�oY[�����%⿄��&(��(����0Z�렿v5Z�����̯��xQ�_'��ʻ��iZ�����T$S����P   P   �^���BH��u���-�ώ���C���S�6[C�~ �1Z�_̘��EG�����J��A�9�1�W˽#��� ;�X@��P   P   .@־ҍ)�uV��Vɿv%���C�nIf��!f�7[C� ���jȿ҃�A�(�4Aվ����=����F&�v�>�ő��P   P   6\��G�soT�K��ϳ��V(�T�oIf���S��(�9�=�����S�u�
�9Ͼ��/��2	��|\w��%���x��P   P   J�Ѿ�&���c'�eu��|���: ��V(���C���C��&(�� �����zt��'�����[nѾ݈;˞Ӿ��Ӿ؉;P   P   T��K2��"�F8�"����|��ѳ�x%�Ҏ���z� C���}����7�L��6�'����)�،3�ǡ)�P   P   xq�K<�]P���G8�gu�M��Yɿ�-�%⿢ɿ�硿��t�r�7����c��<�Nq�n@���5��P   P   S���������L�^P��"��c'�voT�wV���u������Uo���L���[T�;W'��#��c�r�L��ّ����PԿP   P   ��5�տ����M<�M2��&��G�Ս)��BH�uY[��W[�>H���)�DD��*��;�t�<��ˑ��տ���P   P   ��t��1^��&#� 9��4�M�T,�^�����@���ݬ־o�߾E�־/����뫾̰���ﾧ�M��+��#��,^�P   P   �,^��6^�75�S�l��p��՟�N�v���y�\>���C��EC��[=���y�/�v�����|��	��>��4�P   P   #�U�5��:#��i��U��� ��Ġ�8�F�ա'�	2���D�BgM��E�Z2���'�d�F�����d�����?�P   P   �+����,��m���,���+�3A���#5��A������|�Ӌ�$��*���콕B��_�4���d����P   P   ��M�������l-��WN���������4��;ཚ�������Ͻ?	ؽ~KϽ+s��#��̉�^�4�����}��P   P   ������9�%�9�g���B�&���(dF�`\��8$������������kϵ���������!���B��c�F�����P   P   ˰��T,��
�l@�i�
����;b��K�u�*�&���z�����������M���̓������(s���콵�'�,�v�P   P   �뫾��-�� ����N���f߾2��nix�-�0��b�	�ͽ����(��M���jϵ�{KϽ'��U2��y�P   P   *������'��+4�c�<�C�3�&�����e��� =��5OC��B�Fֽ�����������;	ؽ!���E�W=��P   P   ?�־���|,=���b�%y��x��,b���<�
�Xվ� ��&�K��B�	�ͽ��������ϽЋ�=gM�AC��P   P   j�߾w���W��9��;X��OŦ����{ۇ�~�V�Ħ��)޾� ��5OC��b�{����������|���D��C��P   P   ج־�x�t�a�/����繿C'п4п~��������`�Ŧ�Xվ=��.�0���7$���������	2�Y>��P   P   <�����'�W�V���õĿ2�����3c꿐AĿ����V�
�f���oix�*�&�\\���;ཉA��ѡ'���y�P   P   ������9=�?G�����+������3c����|ۇ���<�����2��I�u�$dF���4��#5�2�F�H�v�P   P   Z���oྈ����b��x���Wп������!���6п����,b�'��f߾8b��!�������-A���Ġ�՟�P   P   O,�J"较0��G4��Qy�����Wп-��5��F'пRŦ��x�E�3�N������B����+� �l��P   P   /�M���؇
�r���<��Qy��x�����ŵĿ�繿=X��)y�e�<����h�
�b��ON��,���U��h��P   P   9��D���ڱ9��.�r��G4���b�@G��Y���1����9��Ŧb�+4�� �j@� �9�g-��m���i�S�P   P   �&#�ّ�pv��۱9�ه
��0�����9=�+�W�x�a���W��,=�*��-��
���9����%���:#�35�P   P   �1^�:�5�ڑ�E�����N"�r��������x�w���������S,��������Q�5��6^�P   P   �Ω����aAj��w�Gψ�J|
�����xf��"��&���:��>������[����s
��ǈ��q��:j����P   P   ���������I(,�0����).��Ҵ���l��vV��e�Cv�Zv��e�vZV�?�l�Z�����-�x���,��Ѐ�P   P   �:j�����]j��9,���ǿ>I���Ⱦ�`�4:)�7�)��9���@�59���)�Q)�O�_���Ⱦ��H�k�ǿ�,�P   P   �q��>-��R-�����ݴ�-UI���Ҿ<a���p������� ��� �������N��/�`�Ҿ��H�x��P   P   �ǈ�u>���ο�q���
��*\.�,ɾV�`�ˋ�e���������&K���J��%���r�/�`���Ⱦ��-�P   P   �s
���=���`���`� �=�c�
�sܴ���_�L������_��X�
�Ao�i}�E�$���%��N��O�_�[���P   P   �:��3
�0��e9
�>��iب��l�t|(����3���
�vl���ӝ�E�J�����O)�>�l�P   P   �[��$����aݾ!�����'ݾkP���݌��EU��(�(��+N�#������i}��������)�sZV�P   P   ���� ���?����}�-��O��E���L���Ed���7�v����#�vl�Ao�&K��� �29��e�P   P   ;���6Ӿ�&�bS�^�(�R�(�������1Ҿa����Ht��?�v��,N���
�X�
������ ���@�Vv�P   P   �:��y�㾋4�{�5�xBO�g�X���N�(w5�����y�K$���Ht���7�)���3��_���������9�?v�P   P   #�����ޖ�e�F���m�����͐��tpm�A)F�����y�a����Ed��(������d���n��4�)��e�P   P   
"�� ?Ӿ@:���F�ʚy�2T������*-���y�B)F�����1Ҿ�L���EU�r|(�I��ȋ���1:)��vV�P   P   uf�����	/�� 6���m�$^��>՟���*-��upm�)w5����E���݌��l���_�O�`�5a��`���l�P   P   ����ǰ���J�g�3hO�b���+З�>՟�����ΐ����N���O��iP��eب�mܴ�$ɾ��Ҿ��Ⱦ�Ҵ�P   P   G|
���㾙Tݾ����$)���X�c���%^��3T������i�X�S�(�-��'ݾ8��^�
�#\.�%UI��=I��).�P   P   Dψ���=��
�U��Қ��$)�5hO� �m�̚y���m�zBO�`�(��}����a9
��=��
���ݴ���ǿ+���P   P   �w����@E`�k��U�����g�� 6���F�h�F�}�5�dS���!��,���`��q������9,�D(,�P   P   _Aj�j%-�w�ͿAE`��
��Tݾ�J�
/�C:�����4��&��?澸aݾ3
���`��ο�R-��]j����P   P   ������k%-������=����ʰ�����?Ӿ���}���6Ӿ� ��%���7�㾦�=�p>���>-�������P   P   �d���<���
����.��A��������L�v�v�q�����v;��-�����q���v�Ԧ��j��y=����.�^	���;��P   P   �;��'B�������[V��P��=O���ʾz\t�#�N�]SW�-�d���d��7W��{N�=t��oʾ��N���3V�卵�P   P   `	��ʜ�R��qV�����U�u�=��r���C�*�A���Q�ĦY�-�Q�ӤA�{EC�`.��Ɩ��u�U���3V�P   P   ��.�-�V���V��.�v�⿙�u�����4���D��5;��M�2]���\�- M�);��$D��؋��
���u���P   P   }=��i��L������՘���O�@��1���IF��:��O��f�-�p���f���N���:�+�E��؋�ǖ���N�P   P   m����V�*��������6W�h���ʾb��t;D���:��rP�i7n���������En�<�P���:��$D�a.���oʾP   P   ֦�����	
��7�
�I��R�����s���B�B�:��N��n��Z��؇���j���En���N�);�{EC�?t�P   P   ��v�jk��%���t�̾�̾�}���5���u�߸M�l�@�3LL��*f��р�3z��؇��������f�- M�ҤA��{N�P   P   ��q�༎�茶u&��4�þn�Ջ���6��f\p���U���P�[\�K�o��р��Z�����-�p���\�+�Q��7W�P   P   ,���9ę�����}�о�ྡnྦkоF�q ���ۀ�jc��kX�[\��*f��n�j7n��f�2]�æY���d�P   P   t;��me����ɾj�_��
�e1��,�*�Ⱦh��m_��jc���P�3LL��N��rP��O��M���Q�+�d�P   P   �����h��G�ѾBq�l��2�#��x#�������оh���ۀ���U�l�@�B�:���:��:��5;�)�A�\SW�P   P   s�q�n̙���ɾ;u�	��u�2���:���2��]��+�Ⱦq ��f\p�޸M���B�r;D��IF��D��C�!�N�P   P   I�v�2Ď��������\��Q�2��KC�6C���2�����,�F��6��|�u���s��a���1���4���r��v\t�P   P   ���Lg����V�о�v�g�#�O�:��KC���:��x#�e1��kоԋ���5��M�����ʾ@����7��ʾP   P   ����z�z���)��A����
�h�#�R�2�v�2�3�#��
��n�m��}��B��b�ۉO���u�M�u��=O�P   P   �A���V�%�	�b|̾��þA�ྱv�]����m���_���4�þ�̾
��6W�͘��m�⿿����P�P   P   ��.�`W俨U�����b|̾�)��W�о���<u�Cq�m���оu&��q�̾�7���������.�qV��[V�P   P   �
��!�V������U��&�	�z���𧾻����ɾJ�Ѿ��ɾ����茶#����	
�%���C�����V�O������P   P   �<��y���"�V�bW��V��z�Ng��4Ď�p̙��h��oe��;ę�Ἆ�ik������V�b��(�V�ʜ�%B��P   P   ����i��%���m�;�f���[!�c㧾�j��Z_�0�m�l�u���m��5_�:�j�ѧ��V!�� ����;�v����j��P   P   �j���p����\f�����^��ھ�ⅾ؂e��o���~���~�F�o�?e� ����Dھ�v^�S�����e����P   P   w������1��� 5f�����f����v���y�y��M������,���S���W,���dy��W���q�����]���e�P   P   ��;�%f��5f�q<�)K���z���n�����T���䊾�%���]��#U����ú�����Ғ�������V���P   P   � ��T��r��&K������_������h���x���ڧ�U0��_5ľ�#��a§�k⑾:i��Ӓ���q��v^�P   P   �V!�9�^��d��_x��t_�հ!��ھ����J6����㴬���Ⱦ�ھKھK�Ⱦu���k⑾��� X���DھP   P   ѧ�nyھ����c������ھ���}����Hy�n���P����Ⱦ&>�����E�L�Ⱦa§�ĺ���dy����P   P   <�j��ǅ�Z���ު��ݪ�"�������qKj�:�d�7��Cƚ�F*�پ������Kھ�#����W,��?e�P   P   �5_�OIe���y�&��s�������x��d��D^���n��*��K�n�þ+�پ'>��ھ_5ľ$U��S���E�o�P   P   ��m��o��'�������ȑ�����^���T��wn�5l��}��l��K�G�Ⱦ��ȾV0���]��,�����~�P   P   j�u��~�ד����#����c��<T��w���튾�M}�,#t��}��*��Dƚ�P���䴬��ڧ��%��������~�P   P   /�m���~��㐾�5��G�iȾEȾ6���ܜ���-���M}�5l���n�7��n�����x���䊾�M���o�P   P   �Z_���o�j����;��cľR�پ���q�پ�þܜ���튾�wn��D^�9�d��Hy�I6��g����T��x�y�ׂe�P   P   �j�\e�(1��
��5����پb��r�q�پ6���w���T��d�mKj�z������������s����ⅾP   P   a㧾DÅ�~|y�*���P�����Ⱦ��c�뾼��EȾ<T���^����x�������� �ھ����n����ھP   P   �[!�kPھe��J��/呾נ����Ⱦ��پS�پiȾ�c�������������ھϰ!��_��z���f���^�P   P   c��yw^��u�=���ss��0呾Q���6��dľI�$����ȑ�s���ݪ����k_����!K��������P   P   k�;����<���>���J��*������;���5���󚾈���&��ު��c�Zx��K��l<�5f�Xf�P   P   $�����e��[�=���u�e��|y�)1��k����㐾ؓ���'����y�W�������d��m���5f�.�����P   P   �i������e����|w^�nPھEÅ�\e���o���~��~��o�OIe��ǅ�iyھ3�^�M��!f�����p��P   P    g���<���	����.��>��
�������v�R�q�����:��F����~q���v��������D��a�.�2��f?��P   P   g?��D��˜��V�����V�!��m����ގ�����Av��'k��C������Q��j�+�V��[���V�G���P   P   3��Ͷ�������V�����e���
�ĸ��!��ö�k�ɾ��Ѿӧɾ����ܧ��d����	��U��8�����V�P   P   d�.��_V��tV���.�d��槀��J�4�̾Ii��B#Ѿ�ﾨ��G��n��о����f̾����U�� \�P   P   D��U⿇���͕�?���bCW�0
���̾*ľ���)������3�pz���o�þ�f̾��	�-�V�P   P   ���S<O�#�u���u���O�$�n������G��M����
�N�#���2�;�2���#�ڶ
�������d��j�P   P   ������ʾ�ﾢ����<ﾎ�ʾ�ק��g��ܧ���оw���#�)�:���C��:���#�pz���оܧ�Q��P   P   ��v��*t�bZ���� ���Y���t�_3v�,w���Q�������2���C���C�;�2�3�n�������P   P   �~q�puN�qRC�U?D�
F��D�Q�B�I�M��p�'M��x8ɾ�U�����2�*�:���2����H��ӧɾD���P   P   F���q%W�P�A���:�Rm:��?:�d:�@�@��V��	��9ӣ�^5Ѿ�U������#�O�#�������Ѿ'k��P   P   �:��(�d��~Q�h�L�\�N��P��<N�\L��cP�׃c�4���9ӣ�x8ɾ��w���
�*����l�ɾBv��P   P   ���$�d��Y���\��bf���m�/�m��e���[�yIX�׃c��	��'M���Q����оM�ྷ��C#Ѿö�����P   P   R�q��CW���Q��\�Kp�Ȁ�&������Y�o���[��cP��V��p�,w��ܧ��G��*ľIi���!���ގ�P   P   ��v�}�N�
�A���L���f�hՀ��S���<�������e�\L�?�@�F�M�[3v��g�������̾1�̾ĸ�l���P   P   ����.t�uVC��;���N��n��C���S��&��/�m��<N�d:�M�B��t��ק�h��0
��J�
���P   P   �� {ʾ8���0D���:��qP��n�iՀ�Ȁ���m��P��?:��D��Y����ʾ$�[CW�⧀�b����V�P   P   �>�� O����ߋ��F���:���N���f�Kp��bf�\�N�Qm:�
F�����<ﾍ�O�9���]��������P   P   ��.����u�H���ߋ��0D��;���L��\���\�i�L���:�R?D���������u�ŕ���.���V��V�P   P   �	��x2V�����u���8��vVC�
�A���Q��Y��~Q�P�A�oRC�_Z�����u�����tV����˜�P   P   �<�����y2V��� O�"{ʾ�.t�~�N��CW�$�d�(�d�q%W�ouN��*t���ʾN<O�U⿛_V�˶��D��P   P   �ѩ�2��
>j��s�]ˈ�h}
�����u���.����87������S��G��4ި�5t
�AЈ�"|��Gj�o��P   P   o�����!��B-�D����=�����ڶ�J*��XӾ�����m*Ӿ�輾*����p�k�=�����*-�S��P   P   �Gj�P��_cj�W-�Aο�`��J
�*�ݾ&�澏F�M�!���8�t"�%澸.ݾ;
��?`���Ϳ�*-�P   P   $|��-,��>,�`��kz����`����|m�����'��r6���F���F���5��W���c�������?`����P   P   DЈ�ϳ��ȿ�䴿���d>��X
�f����B)��O��n���y��n�feO�?)�7��d���;
�m�=�P   P   7t
��'.��@I��[I��g.�+�
���㾅�ݾ����2)��
Y�fւ��}��+y��9ʂ���X�?)����.ݾ�p�P   P   7ި������Ⱦ��Ҿ�ɾ$����
�����7,�Z�kO��΂�������엿9ʂ�geO��W��%�+���P   P   G���l���_�~�`�.�`�S�_��bl� �������G�5�H�m�t��������+y���n���5�t"��輾P   P   T��)<V��)�?��Zj�9��2�(�E�U�������Ҿ��V�F�C�y�t�����}����y���F��8�n*ӾP   P   ����ɰe��)��m�Ή��M8�������(�߫d�\���	�W�V�F�H�m��΂�gւ��n���F�"����P   P   97����u�A�8�֐�Cj�&���H	����@�7��t�1����	���H�5�kO��
Y��O�s6�M����P   P   ��uv�Nj@�� �Y����
�Sh
�� ���=?��t�\����Ҿ��Z��2)�B)�(���F�XӾP   P   �.����e�9�� ����,��#�����a���?�7�߫d��������7,澄�������'��K*��P   P   �u���tV���)����(���F����v������ ������(�C�U�~ �������ݾf��{m��*�ݾ�ڶ�P   P   �����l��)�ۗ�����
��f�����#�Sh
�G	����/�(��bl��
����㾃X
�����J
����P   P   g}
�5����_������������
��F��,���
�$���I8��5��L�_����'�
�_>���`��`���=�P   P   [ˈ�]�-�q�Ⱦ�`�$z��������(����Z��Cj�ˉ��Wj�&�`��ɾ�g.����fz��=οD��P   P   �s�z��A�H��Ҿ�`����ۗ����� �� �֐��m�<��w�`���Ҿ�[I��䴿]��W-�B-�P   P   >j��,���ǿB�H�r�Ⱦ�_��)���)�9�Nj@�B�8��)��)���_���Ⱦ�@I�ȿ�>,�[cj� ��P   P   1��bҀ��,� z��^�-�6�����l��tV���e�uv���u�ɰe�'<V��l�����'.�ʳ���-,�O�����P   P   1�t�:3^��##�d2����M�9�"ϯ��	������|�־�߾'�־Ӕ��;ë�����F�*�M��>��7-#��9^�P   P   �9^�>>^�w�5�|���n��MZ辰6���������}�Qq�b��Ye����߾���@��Q���E���5�P   P   8-#�65�]A#�T��1�����9���
�T����-U=���W��a���W�=��t��Pn
���9�v��F��P   P   �>���\�Wt��w���8��e:�\g��4�lk4�_�b�Z����������6?��Ʀb�� 4�2���� �9�R���P   P   -�M�����[���4��(N������
�,�P�<��ry�ŏ��C����Ŀ���an���*y�l�<�2��Pn
�A��P   P   I� ���"��4����\yﾠS��9�@K4��\y����<yп��꿈�꿤`п�����*y�� 4�����P   P   ����q���󹠾�D��lԠ�����୯��߾�z�t�b��w���mп� ���A�v����`пan��Ʀb��t���߾P   P   <ë�wv�)�F�V5��5��F�VFv�8���)����<�o0���������A��A�������6?��=�Ze��P   P   Ӕ��+�y�cg'�0���R"�ۋ����&��x��$��<l��KW�~t��,�Ŀ��꿂 �������Ŀ������W�b��P   P   '�־8��i�1��@��f��7��kP��1���J�վ��:xa�~t�������mп=yпD�������a�Qq�P   P   �߾�-����D�qH�ҹ�������������C�g�����޾���KW�o0���w�����ŏ��Z����W��}�P   P   |�־�:���CM��^�Z�νm���B^���ͽ�r��
L�g���J�վ=l���<�u�b��\y��ry�_�b�-U=����P   P   �����A��6�D��r�J�׽�F��"���ϋ��BLֽ�r�
�C����$��)���z�@K4�P�<�lk4��������P   P   �	���z��2��~�(Ͻ����)���֫�ϋ���ͽ����1��x�8����߾�9�,��4�T��6�P   P   "ϯ�k�v���'����wS���_���4���)��"���B^������gP���&�SFv�ޭ���S辙�
�[g���
�LZ�P   P    9��Ɵ�I�F�rT������g���_������F��m������4��Ջ���F�����Wy����b:���9�l��P   P   ��M���
�����4�������xS��)ϽJ�׽Z�νѹ���f��L"ཽ5�hԠ����#N��8��/������P   P   b2�����B��������4�rT����콠~��r��^�qH��@�+���Q5��D���4��4���w��P��y��P   P   �##�U�<��B��
���I�F���'��2�6�D��CM���D�i�1�ag'�%�F�𹠾�"��[��St�[A#�u�5�P   P   93^���4�U뿉�����Ɵ�k�v��z��A���:���-��8��*�y�wv�o���������~\�45�=>^�P   P   Ⱦ��������q�q����Ѿ�����c־Hu��Cn����`U������վ���=eѾ"���q����D��P   P   E��D��c�տ#Ց���<�;R�c��Kc��)�!PH��W[�TE[�WH�_a)�g�`������r<������տP   P   ����ZԿ���Z䑿��L���yK���'���T��e���~������Ze��<���4T��.'�?���4��L����P   P   �q�;���H��
bq���<����F��48�x,u�����1ɿ�>� ,�ɿ�ߡ�"�t���7�����4��r<�P   P   #��ʠ)�Ȕ3�2�)�����[�-@��%8�����ߎ��N��M8�����#�Œ�OS��������7�?����P   P   ?eѾ�t;�ӾƱӾ��;-�Ѿ�1��^'�[�t�~���C ��m(���C���C�"T(�]( �OS��"�t��.'�`���P   P   ����S������fw��%��"j��S3��m#�@T��롿��cc(��<T�Ւf��0T�#T(�Œ��ߡ��4T�g�P   P   ��վ�b��*k>�����L>�;C����վ�?)�;)��'�ȿv�+�C�Y�f�֒f���C��#�ɿ<��`a)�P   P   ���4��u�:�����˽�f��d:�z��������G��7��2�ῡ��+�C��<T���C���� ,�Ze��WH�P   P   `U��ް��R�>����-���ۨ�԰��<R��I��A����Z��^��2��w�cc(��m(�N8��>⿎���TE[�P   P   ���-���I1l��G�������<Ǭ�����k��9���3���Z��7��(�ȿ��C �O���1ɿ�~���W[�P   P   Cn����l�v�|5�wb��6g�����3���<�U=u��9��A����G�;)���롿~����������e��!PH�P   P   Iu����3jl�5P��ýPW��� h������½�<��k��I������?)�@T�[�t�����x,u���T��)�P   P   �c־�T���=S�Ƒ��μ�ᗇ���_���^������3�����;R�y�����վm#�^'��%8��48���'�Lc�P   P   ����s����K;�w��NN�����)i���_�� h���;Ǭ�Ұ���d:�:C��R3���1��-@��F�yK�c��P   P   ��Ѿ������>�{���7 ������ᗇ�PW��6g������ۨ��f�L>� j��*�Ѿ�[�����:R�P   P   p��8{;����N�q�˽7 ��NN���μ��ýwb������-���˽���%����;�����<���L���<�P   P   �q���)�fӾ�Fw��N�{���w��Ƒ�6P�|5��G�=��������fw�±Ӿ/�)�bq�X䑿!Ց�P   P   �����@W3�fӾ�����>��K;��=S�3jl�l�v�I1l��R�t�:�'k>�����ӾŔ3��H�����a�տP   P   ����8Կ����)�9{;����s����T�������-����ް�4���b���S���t;Ƞ)�;���ZԿD��P   P   �J�� ��Q��z�tG۾ &þ�`ؾd���9!���7�<@��}7��� �dt���׾ʱ¾��ھaf��	Q�_��P   P   _������d�'	.����e��{?,�tx[���@ґ�pđ�p�x[��+�������G����-���d�P   P   �	Q� �`��&Q�.����w��4����N�'e������Կ&���{Կ"J��H ���sN�f���S�V���-�P   P   bf�5s"�f�"�N���'�=���$��c�Q���m!⿴����'���'�Ӷ�����M���c��g$��S�G��P   P   ��ھ�yܾH.��ܾS۾kM�j���}c�r����& ��/5��Pf���z�'f�T�4�N���s@���c�f�����P   P   ʱ¾۟��8���I�������¾��c�N��}��� ���C��^���7��f,���C��ѝC�N����M���sN����P   P   ��׾���`mX��C��X������׾��+�`,����5�U���ص��E��|˵��C��T�4����H ���+�P   P   dt�K[��I(G�����jG��8���Y���Z�*6��2��l f�{+��F���E��f,��'f�Ӷ�"J��w[�P   P   �� ������]�t��Qvؽ�N��t]����� ����>Կ��'�Ǻz�{+���ص��7����z���'��{Կp�P   P   �}7�U-߾g%��8��Ϙ���C��|s�ѵ����޾�7��z���@���'�m f�U���^���Pf���'�&��ođ�P   P   <@�M��4�����(��ǽ$욽a�ƽ�2(�5䑾`��?��z���>Կ2��5���C��/5�����Կ@ґ�P   P   ��7���oܘ�N�6�3ս����qI����ӽ��5��!��`��7���*6����� ��& �m!������P   P   �9!��s߾>�����6���۽������]�'���4ڽ��5�5䑾��޾� ���Z�a,���}��r���Q���'e��tx[�P   P   d��{��Ui��_)���ս�ʉ�Q�L���K�'�����ӽ�2(�ѵ��~����Y���+�c�N��}c��c���N�|?,�P   P   �`ؾ�ş���^�����Ƚn�����^�R�L���]�qI��`�ƽ{s��t]��8����׾~��i���$�4����P   P    &þR����G�Y%���½h4��n����ʉ���������$욽�C���N�gG������¾jM�<��v���e�P   P   sG۾4����X��� �ٽ��½��Ƚ��ս��۽3ս�ǽΘ��Ovؽ���X����S۾�'������P   P   �z���ܾ�H����C���Z%���_)���6�O�6���(�8��s�����C��I��ܾ߬L��.�&	.�P   P   Q�f"����H����X��G���^�Ui��>���pܘ�4���g%����]�H(G�^mX��8��E.�d�"��&Q��d�P   P    ���`�f"���ܾ5��R����ş�{���s߾��M��U-߾���K[�����۟��yܾ4s"��`����P   P   Ms�6�����Ἶ�k��{�¾����?���rE�Yb�X,m��)b��!E��L��.��H>¾H�,��� ��q	�P   P   q	�7�����`�־�P;<5����BQO��
���p���a���M���<���Ǉ���N�e��5z龿�̾b�־����P   P   �侣���徰�־0=پ�� �}�.���y�Q�������_�*?��?�7(��9���y��r.�qu ���ؾc�־P   P   -�������_���Qܼ�tA;\� ��7�������Ͽ���2?L�q�v�p���K�yY�+mϿ�Y��,�6�qu ���̾P   P   I�8���=[��q甾$G�����`�.�������ܿ�N/�*��7X���ڿ�f3��݃�q�.��ܿ�Y���r.�5z�P   P   H>¾Ւ��'�]���]�м��Ƅ¾Ŷ�Tuy�$�Ͽ;/��������c� ��� �9���ƃ��q�.�+mϿ�y�d��P   P   �.��[ ����I��g+��I�C1��DJ��z�N��R���s�!���$��-1�fq��%�9���݃�xY��9����N�P   P   �L����֩\��f�_[���\�Ӂ��x5�񸇿U�U�K��1��!� ��q�fq��� �e3����K�6(��Ǉ�P   P   �!E�������>��%0��W��xL���5澩�D����y���p�����!� �,1�c� ��ڿ�v�p��?��<��P   P   �)b���'���T6�Ͻ�:h�>�5�s���Wd�x�a�������p��1��$�����7X��q�*?��M��P   P   W,m����b�����N�=����½�n����M��U��}p�w�l��y�U�K�!�������*��1?L��_��a��P   P   
Yb�6���}��oL^�t�����2N��gB��4]�����}p�x�a����U��s�;/��N/��������p��P   P   �rE�����+��>v^�]�����Jg��|%��1��4]��U��Wd���D�񸇿�R��$�Ͽ��ܿ��ϿQ����
��P   P   ?����ss��HO��5�AO���'w�B^v�|%��gB���M�r����5�x5�z�N�Tuy�����������y�BQO�P   P   �����0������D7�`c����������'w�Jg��2N���n��>�5�wL��ҁ��CJ��Ŷ�`�.��7�}�.����P   P   z�¾G���֍]��� ��G�sĽ����BO�����������½9h�V����\�B1��ń¾���\� ��� �;5�P   P   �k������wbJ�c2������G�ac���5�^�u��=��Ͻ�#0��^[��I�μ��"G��rA;/=پ�P;P   P   �Ἶ����T^��,�c2��� �E7�HO�?v^�qL^���N��T6�>���f��g+���]�o甾Oܼ���־_�־P   P   ��侞���
~���T^�wbJ�֍]�����ts���+���}��c���(�����֩\���I�%�]�;[��]����徱���P   P   6�� �����������H����0���群��6�������������[ ��Ԓ��7����������6�P   P   <����,��Zy��u�z=����ʾm
���7��Qe�x��|���jヿ��d�%B7��	�r,ʾ@������S2�����P   P   ���� ���(��5 ���8������)�_�n����
ƿF޿+޿R�ſ�Z��dAn��j)�͙����ō���戾P   P   T2��E~�Ud��<���,��²���A��z��4bѿ8��0~0��M>��N0�����п����@� >�1���ō��P   P   �����d���d�ñ������nKJ��Ο�h����>��c���/��W��L.���x>��s���[����I� >�����P   P   @����H_�9DF���_�*����0`A����.���`����������}������6`�ۏ��[����@�͙�P   P   r,ʾ��}��;�� ;�~�S�ʾұ)��K��t���!�`�w��]�#e.�"X.�[;�����6`��s�����j)�P   P   �	�S~��u�K��'��L������
�Xmn��ѿ.�>��ð�VS�B?���P��2?�[;�����x>���пdAn�P   P   %B7�	Ӿ)|w�eD(�A<(��cw���Ҿ=47��R��	���.������QZ.���P���P�"X.�|���K.�����Z��P   P   ��d��g����;�����f;�Vm��{���d�(�ſ�"0�����[x�QZ.�B?�"e.����V���N0�Q�ſP   P   jヿE���0�X��_�h6�8$X� ���S��������ݿ�=���������VS�]������/���M>�+޿P   P   {����+�(�ξ�t�������;�?�s�-
ξ��*�h*����ݿ�"0��.���ð�v�����c��/~0�F޿P   P   w��G0+�s$׾�Ă�C���\۽��ڽ����5���S־��*�����(�ſ	��.�>�!�`��`���>�7��
ƿP   P   �Qe�:���ξ�܂�{�!�@Oҽ$���sѽ|� ��5��-
ξS���d��R���ѿs���-��g��3bѿ���P   P   ��7�~V�et���u�2��P�ҽ%~�����sѽ���?�s� ���z��=47�Xmn��K������Ο��z��^�n�P   P   m
���Ӿ�,��YtY��I�gܽ�E��%~��%�����ڽ�;�7$X�Vm����Ҿ�
�ұ)�`A�mKJ���A���)�P   P   ��ʾ�)����x���<��C�!D��gܽR�ҽBOҽ�\۽���h6��f;��cw�����S�ʾ�0���²���P   P   y=����~�WM�!I)�����C��I�3��|�!�D�����_����@<(��L�~�)������,���8��P   P   u�)`�z�;�� (�"I)���<�[tY��u��܂��Ă��t�1�X��;�eD(��'�� ;���_�m̃�;���5 ��P   P   Yy��nGe�]�F�{�;�WM���x��,��ft����ξt$׾)�ξ��g���)|w�u�K��;�7DF���d�Td���(��P   P   �,��K�~�nGe�)`���~��)����ӾV�:�H0+��+�F��	ӾS~����}��H_���d�E~�� ��P   P   �+����ޗ&�|S�����2Ծ�n�:H�F�z�ٓ���Η�xp���>z�$�G�x���CӾ�����aR�q�%��z�P   P   �z����*���`��h�������p6�p3��F����xۿ1r��Q��p$ۿG:���΁���5����������_�t)�P   P   r�%����kP&�	�`��Z������O��̝�Dk过!���I��Z�(qI�~� �G�翲K��D_N��6�R����_�P   P   �aR�}=��t��
S��:������JX�b箿�{��E[��2���޼��¼�K��P�Z�6�Q[���W��6�����P   P   �����>��I��Z?�)��7}��^�N�@Ԯ�BJ��`��"��,�68�1����X	�����Q[��D_N�����P   P   �CӾdX|� �/� �/���|�̫ӾB!6�I���\�HQ������L*���K���K���)�܅��X	��6��K����5�P   P   w��/E���yU���,���U�)m��,�x���G
�L�Z�����7*��^�z�p��^���)����O�Z�F���΁�P   P   #�G����ւ��qR9��O9�3�����S�G�
>��i� �/���y���K���p�z�p���K�0�K��}� �F:��P   P   �>z�({��㩾��S�8+��kS�,����U�z��ڿ*GI�9����&���K��^���K�58��¼�'qI�n$ۿP   P   wp����+�g˾yt�̽)��)��t���ʾ3G+�{1�������2Z�9���x�6*�K*�,��޼��Z�Q��P   P   �Η���:��`��9��X�/��;�Xj/�Ո���⾉f:��t������*GI�/����������� ���2����I�/r��P   P   ؓ��]�:�S_�.���7� P���{b6�"����뾈f:�{1���ڿi� �K�Z�GQ���`���E[��!��xۿP   P   D�z�-�+�(��.I��N::�������սa����]9�"������2G+�z�	>��F
�\�BJ��{�Ck�D���P   P   :H���B�˾L����f7�� ����ƽ�ƽa���{b6�Ո���ʾ�U�S�G�w���H���?Ԯ�a箿�̝�o3��P   P   �n�W��m��cu�y�0�/��c�ֽ��ƽ��ս��Xj/��t�,������+�A!6�]�N��JX��O��p6�P   P   �2Ծ����)���T���*�d�0��� ������ P��;��)��kS�3��)m��˫Ӿ6}������������P   P   ����}���V�[�:�^,���*�z�0��f7�O::��7�Y�/�ͽ)�8+��O9���U���|�)���:���Z���h��P   P   |S�*@���0�=�-�\�:��T�cu�M���/I��.���9��yt���S�qR9���,��/��Z?��
S��`��`�P   P   ޗ&�� ��! ���0���V��)��n��C�˾*��U_��`�h˾�㩾ւ���yU���/��I��t�jP&��*�P   P   ���y�� �+@��}����Y����.�+�^�:���:���+�){����0E��dX|��>�|=������P   P   p5���C��`����0=�����.&ؾT���M��z��G���U��.ؓ��9��1M����!׾�*��W�;��W���t��P   P   �t���嶽�����1D��A���L��#x:�@B������v��������;7���Մ���9�+*��}i��?	C�b���P   P   �W��:=ͽ]J���D��*��(|�(S�:��%����$���N��s`�ڴN�\�$�~�����GAR�^��[a��?	C�P   P   W�;�؉�}����<�-���k��3\�Ε��ʲ��a��̠�������������x`�t>������l[�^��}i��P   P   �*��{_2������2��������X�R�\����������^^���]�b���9�Y���입�>O�����GAR�**��P   P   !׾��}��5-��^-��)~���׾]):�(	��n������������.�<JQ�o9Q�x�.�Yc��랅�t>������9�P   P   ���_����\��r2���\��ӱ��!�S��.L��`�l8����.�3�c���v�w�c�x�.�X����x`�}�쿊Մ�P   P   /M�\������D�{�D����}�M��G��D�$�퓠��E��BQ�&�v���v�n9Q��9�����[�$�97��P   P   �9���:��豾#b��>9�=�a��Ǳ�� ��%����߿�N�Ai��G���BQ�3�c�;JQ�`������شN��P   P   -ؓ�ɵ0�m�Ӿ9W���x9�pW9��$��S�Ӿ�p0��������#`�Ai���E���.���.��]�����s`����P   P   U���(@��y쾮̑���@��9!�h@�p��y�뾴�?�P�������N�쓠�k8������\^���̠���N����P   P   E���*B@����O�����H�4��MZ��>H��v��������?������߿D�$��`����������a���$�v�P   P   �z����0�C����vfL��u������	���K��v��x���p0��%���G��-L�m�����ɲ�#�����P   P   �M�����]Ծ���A@I�,��{�t�	��>H�p��S�Ӿ� �M�S��'	��[���͕��:��?B��P   P   S��?������ӂ��A�������{｛���MZ�h@��$���Ǳ�|��!�\):�W�R��3\�'S�"x:�P   P   -&ؾ2{��?����Ec��~:��"���-���u�4���9!�pW9�<�a�����ӱ���׾�����k�'|��L��P   P   �����/���]���E��s:��~:��A�B@I�xfL���H���@��x9��>9�z�D���\��)~����,���*���A��P   P   �0=�8�3�Uq.���3���E��Ec��ӂ������Q����̑�:W��$b���D��r2��^-���2���<��D��1D�P   P   _����r���Vq.���]�A�������]ԾE������y�o�Ӿ�豾����\��5-����|��[J������P   P   �C���Tν�r�:�3��/�3{��A�����0�,B@��(@�˵0��:�^�`�����}�z_2�؉�9=ͽ�嶽P   P   ��`�̒����׽��0��c��)�Ҿ�G��F�7�v�Ǐ��\��aj��dQv�F�O����Ѿχ��v�/�y�ս����P   P   µ��4-����ѽ�I5�e"��%�@a4����ê��ӿ���mt�Lӿ�U��x�~�֨3���ﾉB��F4�{�нP   P   z�սz(����ֽ�5��t���8��uK��ʙ�a�߿U"�;%>�zM���=���{�޿mA��\�J�Ţ �=���F4�P   P   v�/����	�k0�,�(�NT�����x$��M�t9���������U����XM�0���$��C:S�Ţ ��B��P   P   ·���H*�����*�������LK�����
��Ys�eY�������������A�r�۬��$��[�J����P   P   ��Ѿ�.x��R)��)�y�x��XҾ�4������
�vAs��S��i��/�=��=��~�����A�r�/��mA��ը3�P   P   N��酮���Z�&�1���Z��Ʈ����E�3G߿��M�X:������O���a�}�O��~�����XM�z�޿w�~�P   P    F�������E���E�����>�5F�p��.��������W�=�$b���a��=���T������U��P   P   bQv��i��7���Yd�Z<=��Dd�^#���Z�3<v�;ӿ'�=������W�=���O�.�=����������=��LӿP   P   _j����+�>AѾX烾k�@��d@�μ��/�о![+��@��
/�=M��������h��������zM�jt�P   P   \��R3:�L,�̓�4K���-��J��x��{��n�9�4��
/�&�=����V:���S��cY��r9��9%>����P   P   ŏ��lL:����I����U�j\'�A*'��^U��Μ�W�n�9��@��;ӿ.����M�tAs��Ys���M�S"��ӿP   P   5�v��+�s�g���Z��&�0K��=&�A�Y��Μ�{��![+�2<v�p��2G߿�
��w$�^�߿�ê�P   P   �F����5�Ѿ���ZV�u�&�V��2���=&��^U��x��/�о�Z�5F��E��������������ʙ���P   P   �G�t�᰾�e����K���'����W��0K�B*'��J�μ��]#���>����4��LK�MT��uK�>a4�P   P   '�Ҿ�h��������e�:�A��.���'�v�&��&�j\'���-��d@��Dd�����Ʈ��XҾ����(��8�"�P   P   �c����y��!\��G��p>�;�A���K��ZV��Z���U�5K�l�@�Z<=���E���Z�x�x���+�t��d"��P   P   ��0�Ø+���*��2��G���e��e�� ��g���I��̓�Y烾�Yd���E�&�1��)��*�k0��5��I5�P   P   ��׽�{�
����*��!\�����᰾7�Ѿs龿�N,�@AѾ�7������Z��R)�����	齽�ֽ��ѽP   P   ˒��V���{�Ę+���y��h��w�����+�nL:�T3:���+��i���ꅮ��.x��H*���y(��3-��P   P   9�4��tg�����%#�8n��mKþ�8	��4�M�^��;~��넿�}��^��s4�T���I¾�����!����Զe�P   P   նe�[�f��h����&������޾��$�ղf�O����a���fο�IοK���Y����e��H$���ݾu8���T%�~���P   P   ������p	���Y&�����sz�Zg9�����!ÿ�\�����3*������¿v���8��Z�w0���T%�P   P   �!�-JӽH�ӽ��"��⌾�]�n�@�����H�濏}*��i�1������h��
*��<�nz���5@��Z�u8��P   P   ������K���K����h]޾-D9��򖿭���8F�U������R������� ����E�c`��nz���8���ݾP   P   �I¾x7g�p�u2���g���¾��$�Ol����濆'F�nf��8M���O��@�~ ��2����E��<�v���H$�P   P   T��PD����L��'�i(M�����>���Sf�	�¿�T*�?��PB���z%�?�5��f%�} �����
*��¿��e�P   P   �s4���׾\V��ɾ;�d�;��k����׾�4�Hx�� /���h����sL�b�5�?�5��@������h����Y��P   P   �^�v��󭥾7�[��T8�:�[�����j��Ӏ^�����z�
������sL��z%��O�O�������I��P   P   �}�����*žƀ�k�B��B�4�����ľ&���}�vο*�
������NB��6M������/����3*��IοP   P   �넿O�*�,ܾ9:��%)V��=���U�X둾��۾,�*�d���vο�z���h�?��lf��U���i�����fοP   P   �;~���*��侯֜��h��E���D��g��_����,�*��}�����.��T*��'F��8F��}*��\��a��P   P   J�^����^ܾ��<p��=M��QC�0�L�fo��_����۾%��Ҁ^�Hx���¿��濪��F���!ÿM���P   P   �4�+[�A�ž���H�h�]rM���D�ҕD�0�L��g�X둾��ľj���4��Sf�Nl����~������Ҳf�P   P   �8	���ؾ�P��2A����V�8�E�z�C���D��QC���D���U�4���������׾>����$�,D9�l�@�Xg9���$�P   P   kKþV����6�\���C��>�8�E�]rM��=M��E��=��B�9�[��k��������¾f]޾�]�pz�޾P   P   7n����h�NN��=��}9���C���V�I�h��<p��h�%)V�l�B��T8�c�;�h(M���g�����⌾�������P   P   �%#�)$�sG�?M(��=�8�\�4A�����󜾰֜�::��ƀ�8�[�ɾ;��'�t2��K���"��Y&���&�P   P   ���q:ս�%��tG�NN����P��C�ž ^ܾ��.ܾ�*ž����]V����L�o�J��E�ӽn	���h��P   P   �tg�"H��s:ս+$���h�Y����ؾ-[������*�Q�*����w����׾QD��x7g���,Jӽ���Y�f�P   P   ���	?��k�����d�IЪ�����\�>��X��ea��W�F>���� ��䩾�Bc��O�
ģ�X]=�P   P   Y]=�E>�����A���x���¾#��±D�+`~��瘿G����k��^�����}��D�3*�\�����v�����Z��P   P   ģ��&v�趤�]���3�ܲо� ��yh��E����Ͽ�����0�����[KϿfԟ���g��Z��Ͼ��}����P   P   �O�����0;�����w�>�о�X&���}�����Gr���+���G��G���+�f"����V�|�7�%��Ͼ��v�P   P   �Bc��b	�5ٽ��	�[-d�B�¾��,�}�d�Ŀ���ԖX�4@��4���&���,X�1L��CĿV�|��Z�[���P   P   䩾JAJ��y	�w�	�Q�J��d������Dh�K������rk�f���2�����A��Mk�1L������g�2*�P   P   ���R3����3�V���84�{x��A��gD�G���X��|X������������a��@���,X�f"�eԟ��D�P   P   ���D���vk��)��))��k�gp��E��n�}��xϿ�+��0��m/��e���������$����+�YKϿ��}�P   P   �E>���쾘����M��O0�b�M�����w��EH>���� ����}G�	���m/�����2��2����G�����]���P   P   �W��U
������{�CK��$K�&{�GI��(4
��W��O����}G��0�����d��2@����G��0��k��P   P   �ea�n���˾/���'s�3�c�@�r�7ؓ��˾#���a��O�� ����+��|X�rk�іX���+�����E���P   P   �X����+Ծ�,�������g��2E���������6�Ӿ"���W�����xϿ�X�������Er��Ͽ�瘿P   P   Y�>���
���˾H��ܚ���1���e��M擾��������˾'4
�EH>�m�}�F��J���b�Ŀ�����E��'`~�P   P   ���������.|��1��WP���z���R��M擾���6ؓ�FI��u��E��gD��Dh�)�}���}��yh���D�P   P   ���	��,��2�|���s�滅�%����z���e��1E��>�r�${�����ep��?��������X&�� �!��P   P   FЪ�����I�l���N��>L���d�滅�WP���1���g��1�c��$K�a�M��k�zx���d��@�¾;�оٲо��¾P   P   �d�E�K�H5�NJ*��i1��>L���s�1��ܚ�������'s�CK��O0��))��84�O�J�X-d���w��3��x�P   P   ��Ԝ
�ϩ
�3��OJ*���N�4�|�/|��H���,��/����{��M��)�U��v�	���	��[��>��P   P   �k��\���� ۽Щ
�	H5�L�l�,��������˾�+Ծ�˾��������vk���3��y	�3ٽ-;��嶤�����P   P   �	?��mx�]���՜
�H�K������	������
���p���U
����D��S3��JAJ��b	������&v�E>�P   P   ���+�c~���E�:��P����þ����@��{�/���6�.h/��6������þ����i9��d�?Z{�|��P   P   |���h��u�[n�v�K�������龚:�*�J�}�p��c��QS��O5p��oJ������辎����J��\齌&s�P   P   @Z{�`"5�9}���cYR�{i��s����:�u({�(��g���|c��ff���ȝ��z��.:��l�΅��}Q��\�P   P   �d�Rċ�#4����{�K��T�����K�0��-�������R	�/B	������������aJ�g��΅���J�P   P   �i9�6ڽЗ����ڽ>:�jW�������J�� ��ڱؿ����5�8IC��4�ޜ��8ؿ�����aJ��l�����P   P   ����#�06ڽ}�ڽxv$�����s��M�:��
��ڥؿQ%���S��2z�z��bS�����8ؿ�����.:����P   P   �þ�Kj�Q����ｼ����j���þ����z�z���!���S�z����ĕ�u����bS�ޜ� ����z����P   P   ����6��SI�;�� ���0I��1�����@�J��읿��5��0z��ȕ��ĕ�}z��4�����ȝ��oJ�P   P   �6��
Ⱦ�-���D��z/��D�$��dȾ�9��?p�tl���C	�&HC��0z�y����2z�5IC�.B	�df��L5p�P   P   ,h/����ͼ������Al�il�?Z���s���n뾉H/�B��\L���C	��5�
�S���S��5��R	�yc��PS��P   P   ��6��C �����,�������:��H��I@��T�� �t�6�B��tl���� ��P%�������d����c��P   P   y�/��T �M�ʾ����ȾS0ؾ��׾�Ǿ�h��2ʾ~ ��H/��?p��읿x���إؿرؿ*���%��y�p�P   P   >��$����-5��h�ؾ: �٦	�����B�׾�h��T���n��9�>�J���z��
��� ��.��r({�'�J�P   P   ������Ⱦ� ��.���[Ⱦ�O �j����������ǾH@���s��cȾ�����K�:���J��K�}�:��:�P   P   ��þw���N����������ؾM�	�j��צ	���׾	H��=Z��"���1����þp�龢����q�����P   P   �P��j�k��9J�`�E�rAm��ˡ��ؾ�O �: �P0ؾ:��el�ߣD��0I���j�����hW���T��xi������P   P   A�:��@%��������0�sAm������[Ⱦf�ؾ�Ⱦ�����Al��z/������vv$��=:�w�K�_YR�r�K�P   P   �佬<ܽ4YܽO�����b�E���.��-5�����+�������D�:�����z�ڽ��ڽ����Vn�P   P   c~�lr���Y��6Yܽ����9J�P���� �����N�ʾ����ͼ���-��SI�Q��/6ڽΗ��!4��4}��u�P   P   *�97�mr���<ܽ�@%�n�k�z�����Ⱦ(��T ��C ���뾏
Ⱦ7���Kj��#�6ڽQċ�^"5��h�P   P   �#���q��-�>�����
��V��	����Ǿ4u���F
��!�F$
�]��'[ǾyW��;&U�'�	�2���w~��Ol�P   P   �Ol��Lo�Jc��ǧ�����w�Qٴ��D������6�{�E��E�|�5�����p��k��?�u�"w�����'.�P   P   w~�d���8������P�]`����ʾ�.�u�<�-�h�rل�����������h��<���w	ʾ����*�����P   P   2���#T.�N/�Y韽	p��O���ӾL�	�V�}���Z�������8���Պ��O���7V�����8Ҿ���!w�P   P   '�	��W���G[���� i
�/�v���ʾB��f`�~���{�ſ���P����n��NſQ����_����v	ʾ>�u�P   P   :&U�{񽚕���ޘ��\���U�ז����h�V�ɖ��Y�п�����s����I�пQ���7V���j��P   P   xW��!5�V�nලگ���5������A�<�������ſ���i� ��,�
� �����NſO���<��p��P   P   %[Ǿ
@~�Q�)�[�DZ�1�)��k~�b�Ǿ#��V�h�d���g�鿒��,���,�r��n�ӊ����h����P   P   Z���J��u�`�M�	C�>SM�Ӿt��-�����}�5�������U�����h� ���M���6�������z�5�P   P   E$
�r�Ⱦ��������hݟ�p����M��	,���wȾ_
�1xE��늿����f����������鿺��������E�P   P   �!���ݾ�qǾ��׾6r���o�����׾װƾ��ܾa��1xE���c�����ſW�пy�ſX���pل�x�E�P   P   �F
�+�ݾ?վ�H �D#(��H�V�H���'��d��oNԾ��ܾ^
�|�5�T�h�����ǖ��|���{���*�h��6�P   P   0u���"ɾ�Ǿ�V �$;��!|�����z�{�VZ:��d��ְƾ�wȾ���"��?�<�e�V��f`��V�q�<����P   P   ��Ǿ���������/ؾ�N(��J|�o���G���y�{���'��׾,���-��`�Ǿ������B�L��.��D��P   P   �	��p\��u��������%SI��׌�n������R�H�����M��Ͼt��k~�묗�Ԗ����ʾ�Ӿ��ʾMٴ�P   P   �V��M6�k�*���N�$n�����$SI��J|��!|�z�H��o�l���9SM�-�)�݅5���U�+�v��O��[`���w�P   P   ��
�E��#Y��O��D�$n�������N(�!;�@#(�/r��dݟ�	C�AZ�կ⽔\��h
�p��P����P   P   :���D���n��ʮ���O���N�����/ؾ�V ��H ���׾����[�M�[�jල�ޘ����U韽�����ǧ�P   P   �-��D1�mX^��n��'Y�n�*� �u������Ǿ?վqǾ����u�O�)��U⽘����G[�I/�3�Ec�P   P   ��q�"dļ�D1�D��K���M6�u\������"ɾ-�ݾ��ݾs�Ⱦ�J��
@~�!5�{�W��!T.�_����Lo�P   P   �Q<�u�;T>��p/�����W��v�]��R���~��:�־�����־���ӕ�`�\����񔱽G/,��&5����;P   P   ���;��;݅1�V=���˽�,.��ق��G�����*�\c��R�����}�Ӥ��x2��v�,���ɽ�D:���)�P   P   �&5�]��9i�:�o�<��bս�=����о����k&���;�ױC�x�;�5$&��W��о����Ѯ<��tӽ�D:�P   P   H/,���g��j��).�^˽�=��虾e����d�D�̈h�ԡ}�
�}�sGh�WDD�j'���ᾩ7��Ѯ<���ɽP   P   񔱽��+����_̲�M�-��{����⾵4!�
�V�ET��������y���5*���5V�� ��������u�,�P   P   ���&���,�>'-������M�c���<�оz���V�:Ë��!��W:���.����������5V�j'��оw2��P   P   _�\��V��ܣ�Į��Q������U]��������D��M��q����ſp�п��ſ���4*��VDD��W�Ҥ��P   P   �ӕ�rKI������B���?���GI����L&��rh�����;���пp�п�.��x���qGh�4$&��}�P   P   ���ь��|u�ys�،v��r�(�t�����q��A����;�X�}������;����ſU:������}�v�;����P   P   ��־l��D�����Ӿ��[�;Ӿo봾�ܱ�B־J=�ߤC�W�}����p���!�����С}�ԱC��R�P   P   ����ɾ���p��-R���h��xQ�����`辀ɾ"]�J=��;��rh��M��8Ë�CT��Ɉh�}�;�Zc�P   P   8�־�ɾ~�����F�ﭖ��%���便��|�E��h��ɾB־A��L&���D���V��V�a�D��k&��*�P   P   �~��l���7����F��媿�C��e�l���� ��{�E��`��ܱ�o�����~��x��4!������}�P   P   �R��-���������Ӗ��l��JB!��!�j���}�����k봾���9�о���a�⾂�о�G��P   P   q�]�(.J� ?v�jBԾ�pR�ք��1X�IB!�b��便�xQ�4Ӿ!�t��GI��U]�a����{���虾앓��ق�P   P   R���K����4
t��l�7ki�Մ���l���C���%���h�[���r�:������M�I�-��=��=��,.�P   P   ��������l������l�w��l��pR�Ӗ��媿ꭖ�%R���Όv�7���K������Y̲�^˽�bս��˽P   P   �p/�-!�-�/�E=�����4
t�hBԾ�����F���F�j����Ӿps��������6'-�
��).�f�<��U=�P   P   	T>���q��̿�1�/�o������?v�����4��y������?����|u����ܣ��,�"�����j�U�:�Ʌ1�P   P   �u�;�)���q�3!������K�,.J�-��m����ɾ�ɾl���ь�qKI��V�%��	��~�g����9/��;P   P   O�	=\ �<O�|<a��P/����+���Z��ˎ���w�����􆎾 /Z�N��a���,� n����<��<P   P   ��<��<ۀ<�:7�8sS��<׽��-�)�v��V��>缾9�;��;K���Z�F�u���,��Lս"P��-�� �<P   P   ��< w�<�<��5�c�u&���E��C��/������V�d��8;�({�r�����x�D��/�%�_��-�P   P   n����d<�b<���W�R����,5O���6վ������*�^�*��w��}��Ծ!����N��/�"P�P   P   �,��b��Au�;wA���.���ֽ
�E������޾A���3�JgJ���R�zHJ��2��R��.޾ ���w�D��LսP   P   �a��z��(VV��W�����U��@p-�^'��LmվD��G�:�:]�� q�\�p�u�\�0�:��R��Ծ�����,�P   P   N�_Ȳ�N�e�W?��f��������^v�|ϼ�����2�m]�"7|�f僿�!|�u�\��2��}�r��D�u�P   P    /Z�	�!�ę�[t��O��G��j!�.1Z����t��ט�>eJ��q��胿f僿[�p�yHJ��w�&{�Y�P   P   􆎾wj{����Ӝ��ޥ�B4��W�����z��K��j���&D��*�fS��q�!7|�� q���R�\�*�6;�I���P   P   ���n���۾���K�7�`�7�D��Yھ�����~���};��*�=eJ�k]�8]�HgJ��*�b����;P   P   w����Ǿk���/r�<����G¿�5��	�p�����Yƾ����};&D�֘���2�E�:��3�����V�6�;P   P   ����Ǿr�&�))������A%��%������,��
p%��Yƾ�~��h���r����B��?���� ��;缾P   P   �ˎ�I���׾�Q6��3����X�`Jx��ZX�t���,����������K�����zϼ�Imվ��޾2վ+����V��P   P   ��Z��{�m�۾�lr��(��|Y�0o��J���ZX������p��Yھ��z�*1Z��^v�['��������C��"�v�P   P    +��X"�Yi��/����ǔ%���x�/o��\Jx��%��5��yD�R����j!�~��<p-��E�'5O��E�~�-�P   P   ���BK���J����f|8�9�¿Ɣ%�yY�|�X�A%��G¿X�7�;4���G�����U����ֽ���m&ｅ<׽P   P   P/�����h��B�����e|8�����(��.������4���B�7��ݥ��O�tf�����.�L�R�c�,sS�P   P   D���-Ż<V`��B��B����/��lr�L6��")���/r����˜��Rt�W?���W�;A��m����5��:7�P   P   _�|<K�\<$��;GV`��h��J�Xi��i�۾Ӿ�l�&�e����۾������@�e�
VV�ju�;%�b<�<'ۀ<P   P   _ �<���<B�\<!.Ż���HK���X"��{�H�����Ǿ�Ǿ�n��qj{��!�[Ȳ�u���b����d<%w�<��<P   P   �Y=�TL=��#=�}�<�����	,��\��˸��\[��Ć�&j��^���<�Z��,����c)���j���<k%=�M=P   P   �M=\�L=  $=ׁ�<� �-�K��ʽ��U��ہ��Q���A������nT� R�3Ƚ��H��c��<�f%=P   P   k%=c�?=V�$=��<�O��sm��(��4��v��◾���1$���ͫ�_���`u�Q4�;k罀Zj�*VE�b��<P   P   ��<��=�{=��<���s<m�=���x�F�m���v���Ͼڞ����}Ͼ���[����E�@��Zj��P   P   ��j��<�=ye�<�⁻�QK�`��4�F��ؑ�&_��Xz��j�خ	��U��+�0����h���E�:k罤�H�P   P   �c)���ĻX�,<�+<�|ʻ8�*�j�ɽ޴4�fb��F[������Y"�����R��y��0���Z���P4�2ȽP   P   ���c�ɜ!�x��d!�ȋc��g�������u��i��w�E#�v�"�Q�)���"�R��+뾫��`u�R�P   P   �,�����eI����t�> ����1�T�j×��Ͼm��%�ζ)�Q�)����U��}Ͼ]����nT�P   P   ?�Z�sm�X����LžF�ؾްľ�����l�dAZ�q���bث���ྖ�	��%�u�"���֮	����ͫ����P   P   `���A���^���=L��؀�S���(HK����7P�������������m�D#�W"��j�֞�/$���A��P   P   'j��(�о�7?�G᩿.��{��}j���ܨ�ȵ=�i�ξê����aث��Ͼw뾖���Uz��Ͼ����Q��P   P   �Ć���о�FW�iݿW:�q�s�\�s���9�O�ۿa{U�g�ξ���o���h×��i��D[��#_���v��}◾�ہ�P   P   �\[�\����I?�`ݿ�U�Ey���
��X����T�M�ۿŵ=�3P��`AZ�-�T���u�db���ؑ�m���v��U�P   P   ȸ�]�m�B����Ն:�d����T��3��W����9��ܨ�����l�������ڴ4�/�F�r�F��4��P   P   �\����?Κ���L������et�YN���T���
��U�s�uj��HK�����8 ��g��c�ɽX��4����(��ʽP   P   �	,���e������ž7;���N��et�a���Ay��h�s�u��M���Ұľ�t���c�+�*��QK�e<m��sm��K�P   P   ?�����ֻ��#���)�پ6;������ц:��U�W:��-���؀�8�ؾw��d!��|ʻ7⁻����O�� �P   P   �}�<C�<��$<d������ž��L����Wݿ_ݿ=᩿�=L�vLžXI��w��+<�e�<��<��<健<P   P   ��#=ZT=m =��$<��#����=Κ�?��I?��FW��7?�V��N�������!���,<�=�{=Z�$=$ $=P   P   �TL=C�>=XT=9�<�ֻ��e���[�m�Y�����о �о:���sm���
�c���Ļ�<��=e�?=^�L=P   P   ��=�L�=Z�u=��@=���<���\�J�Rؽ:**���\�X5p��i\���)���׽��H�%��g�<�}B=�w=ǚ�=P   P   ǚ�=�o�=J�u=(;=r��<Fyƻ�1��˰�`���!,���B�0�B���+�p(�Eů�^/�%����<ν<=��v=P   P   �w=��=�Tv=[W;=k.�<�X4��VS���ƽ���\�<��Y���c��WY��<��;��ŽڠP���*�,�<ν<=P   P   �}B=3�q=�Vq=�qA=�P�<�3�+e�C�ݽ�T'���[�뜂�V����덾�o��Nm[���&�iqܽ�b���*����<P   P   g�<9�9=
�R=�R9=��<B�»�S���ݽ��/��,q��Ҕ� ������� �������p��R/�hqܽ٠P�,�P   P   R���ْ<���<LP�<��<Bi��_�0��ƽ�H'��)q�����
���t�ƾQ�ƾpY��:y���p���&��Ž^/�P   P   ��H�w��oQ伬7�TU��q��I��4��Y����[��Ӕ�y���5�Ͼ�Gؾ��ϾpY������Lm[��;�Fů�P   P   ��׽��彃m�#{(��0(�C��$����ֽ�$��R<�=���s(���ƾ�Qؾ�GؾO�ƾ� ���o���<�p(�P   P   ��)�C�c����	��)� ���V���Bb�>�(���+��]Y���P���ƾ4�Ͼr�ƾ�����덾�WY���+�P   P   �i\�ڳ�����]2u�uV�����Z�s��u��?����Z�6B�f�c� ��r(��w������ ��S�����c�0�B�P   P   _5p�e=ؾ�_��*Ͽ�f�n/�����Ϳ�(]��E־_wn�5B��]Y�<����Ӕ������Ҕ�蜂��Y���B�P   P   ��\� Fؾ0�|�K)��3f��R����u:e�R<��]z��E־��Z���+��R<���[��)q��,q���[�W�<��!,�P   P   :**��ͮ�@_�<5����[���,����H��3=��Q<��(]��?��:�(��$�U���H'���/��T'����]��P   P   Rؽ�4d�+���_Ͽ�pf�۶�����������H��q:e��Ϳ�u�Bb���ֽ�4���ƽ��ݽ:�ݽ��ƽ�˰�P   P   R�J�ҫ��?���u�}������30������*��������O�s�M����但I�R�0�yS�+e�sVS��1�P   P   ³��ܓ������wѝ�*�/�����ض��W����R��f/������7���q��h���»��3��X4��xƻP   P   ���<�x�<��$>)��8�vѝ�z���pf�����3f��f�kV�� � �y0(�U�8��<�<�P�<}.�<���<P   P   �@=$d8=���<+-�#>)����u��_Ͽ75�D)��*ϿL2u����{(�q7�hP�<�R9=�qA=aW;=(;=P   P   ]�u=B{p=7}Q=���<�缆���?��&��6_�"�|��_�������um�9Q伞��<�R=�Vq=�Tv=M�u=P   P   �L�=Z��=@{p= d8=�x�<��ҫ��4d��ͮ��EؾZ=ؾг��5�c����d���ْ<>�9=6�q=��=�o�=P   P   �'�=w��=h��=mЃ=
:C=���<dX�����x��E&3�c3F�3���^�������Ln�<�D=�h�=�'�=�1�=P   P   �1�=��=Fޗ=2�=��D=5y�<E�Q�j������ؽ<=�����6ؽ�򖽰���8����<�CF=��=�@�=P   P   �'�=r�=�ߗ=��=��@=��<�Ͽ�y< ��Օ�L�ӽ V��*w�D���Lӽ����L�&M���?�<�LB=��=P   P   �h�=�ϔ=ѭ�=&�=V�D=	��<U]��/:��⬽j���XS��((��(�������۫�*8�Q� ��?�<�CF=P   P   �D=5�w=���=EFw=�C=8$�<�X��#:�e��'	��/�%J��SS���I���/����궽)8�'M�����<P   P   =n�<�W=�#=p�"=!=O�<�yH����Vլ��'	��"9�Z�^�?Ds�P,s�Rh^���8����۫��L�%8�P   P   ����?i����cj�������ff��7��v	�����������/���^�
�~��9����~�Rh^���/����������P   P   i���
��-�	�PI)� �(�������˒������ԎӽR��.J��\s�FB���9��N,s���I����Lӽ��P   P   ���^R��@���9��6�mh�	.����P�/���i׽�����5(�Q|S��\s�	�~�<Ds��SS��(�A��6ؽP   P   3��ͦ�#� f}�H��^��� |�c��qE���1�j����T��5(��.J���^�W�^�!J��((�(w����P   P   k3F��Ѿ��c��9ֿ����`5�Jr�t�Կ�a��Ͼ�bD�h�������R���/��"9���/�TS��U��<=��P   P   K&3�1#Ѿ�����Ln�Ni��3���Gm�`�
�����Ͼ�1��i׽ώӽ�����'	��'	�b���E�ӽ�ؽP   P   z��,ᦾ��c�����m�������������_�
��a�lE��*����������Oլ�^𷽓⬽�Օ�����P   P   ���юR�S/�'rֿ��n��������������Gm�m�Կ]����P�����i	����:�/:�k< �^�P   P   WX��ؑ��́����}�SG����6������ ���	3��Cr�	 |��-��򁿽q7��$yH�HX��%]��Ͽ���Q�P   P   ���<n�D�	�����ɣ�46� ����������Hi���`5�T���\h�y���ff�(O�<M$�<��<��<Iy�<P   P   :C=h%=�����)����ɣ�PG���n��m��Ln����H���6���(�L���!=�C=^�D=��@=�D=P   P   oЃ=Оv=3�!=˻���)������}� rֿ������9ֿf}��9�>I)�!j����"=MFw=)�=��=4�=P   P   i��=:a�=(��=2�!=����B�	�Ɂ��M/���c������c���@���	�G���#=���=ӭ�=�ߗ=Gޗ=P   P   x��=P��=9a�=͞v=c%=n�Ց��ˎR�%ᦾ%#Ѿ�Ѿ�ͦ��^R����i?i��W=;�w=�ϔ=s�=��=P   P   ���=_��=h(�=+��=�@w=&�=@;0�0��`��Z����m���5���70�i�N;.�=}5x=��=�w�=߮=P   P   ߮=�Ʈ=���=ۘ=��=y<=d�<:���C����z��#��K��bz���[����)�<�==ɂ�=�K�=���=P   P   �w�=_�=�A�=��=w��=ܤ<=���<��9��μYtE�c���S���l���;�D��w̼�r:w�<�>=44�=�K�=P   P   ��=!�=��=n̗=��=±<=���<-h�;���e�����]d��B���Y����c� �����)��<�>=Ȃ�=P   P   x5x=�5�=>7�=��=�w=L�<=f6�<$����F��P���"Xݽ�꽛ݽhl���K���}����u�<�==P   P   %�=N�5=�>=�>=4�5=%V=��<I4�9��������Ž����g
��T
��/���eĽ�K�����r:x)�<P   P   u�N;��\�v���Y�)9���(��U;	����μ�d�;������T��"�L2��/��fl����c��w̼����P   P   �70�e����1�-��������$���L.��Z�X�D�XÛ�Qݽ=~
��1��"��T
��ݽ�Y��;�D�
��P   P   �5����3��(���վgJ�aԾ/���J2�u2��P�x������|���a�<~
�T��g
���B��k���bz�P   P   v���b���q��}`�n䏿����?c_�w^
����s
�
㜽`����|��Oݽ�������XݽXd��Q���O��P   P   ������3I�W����
�1��E
�wY��fzG��/��$Q�	㜽����UÛ�7���ŽJ�������_����#��P   P   `��:	����c������N��K����I�M�9���a��/��
s
�G�x�P�D���d����@��e�OtE���z�P   P   �`��Kp���DI�3��~�l�ꑯ�f\��1,����k�9�bzG����l2���Z��μw���v�"�����μ>��P   P   1�0��4��������PO����@]���=��0,��D�M�qY��r^
��J2��L.������9�9v��ug����9����P   P   G@;�����]����`�� �E�������>]��c\�����E
�4c_��.���$�� U;6��<z6�<���<���<u�<P   P   ,�=������b�վV�����D������呯��K��)������`Ծh��ۻ(�2V=U�<=ʱ<=�<=y<=P   P   �@w=��4=������V?�V��� �JO�t�l���N���
�c䏿TJ����8�C�5=�w=��=z��=��=P   P   -��=�ڋ=Ze==�C^�ߊ�_�վ��`�����'��~��J����}`��վ��Y��>=��=q̗=��=ۘ=P   P   i(�=.Ѣ=}�=Ye==�������]������DI��c��3I��q��(���1�����>=B7�=��=�A�=���=P   P   _��=`�=.Ѣ=�ڋ=��4=��������4�Dp��/	��z���b����3�O�����\�[�5=�5�="�=`�=�Ʈ=P   P   �-�=�p�=|�=�͜=��=�9=ƽ�<t���Ӌ��0�н����{н1v���6��ȁ<��:=�h�=��=��=���=P   P   ���=_{�=%x�=���=ύ=V�e=@Y=�|z<�'�j ��S6�)<6�V �D$��}<�=��f=�0�=�=���=P   P   ��=1Ǭ=L��=���=]��=��l=-=���<��;��W��Ҽ4m��@]Ҽ�IU�¢�;���<� .=��m=K�=�=P   P   ��=K(�=3�=�ڜ=�ԍ=�l=ݺ-=l�<YX�;x�m�A���v��C�����j� J�;?n�<��.=��m=�0�=P   P   �h�=Mڎ=ڤ�=���=�.�= �e=d-=��<b'3;a,���Q�r~K�o]�zK�O}������F;?n�<� .=��f=P   P   z�:=�7D=IxD=�D=
=D=�d:=.�=d�<�q�;6A��h'��Kn�v���Ї��:�m�+ &����!J�;���<�=P   P   �ǁ<$�<�ۺ�5ûn�Ⱥ��<迂< �|<�4�;��m�>p�?kn��8��㟽3��9�m�M}��j����;�}<P   P   �6���a��뿽d<�����������_�˼��{���U����K��̊�4���㟽·��vK�|���IU�l$�P   P   @v��-����u�3d���x���ת�/lt��?��Ɔ��Y����Ѽ��k�]��̊��8��t���o]��C�@]Ҽb �P   P   
|н@Uh���ܾ�`.�/�\��{\���-��ھ� f��νg;4��|�����K�9kn��Kn�j~K��v�0m��3<6�P   P   ��콑
��ε�g���U�ο�����Ϳ\ی�im�C������d;4���Ѽ��8p�`'�xQ�0��	�Ҽ�S6�P   P   <�нI���d0��G��ӎ�*F���E�������5�.�B����ν�Y����U���m�&A��O,��R�m���W�j �P   P   ڋ��ech����<X��{�-�䎁�����;���-����fm�� f��Ɔ��{��4�;;r�;�'3;�X�;=�;�'�P   P   {������"�ܾ�ԍ�K����p������;�����Wی��ھ�?��ʼ�,�|<v�<�<~�<���<}z<P   P   ʽ�<��a�b@v�r�.��Ͽ͖F�@��n��������E���Ϳ��-� lt��_���<8�=l-=�-="-=GY=P   P   �9=��<zQ��Kū�)z]�$��˖F�ꦁ������)F�����{\��ת�����S�<�d:=�e=�l=��l=\�e=P   P   ��=��C= !��D,��'z]��ϿF��t�-�ˎ�H�ο �\��x��l����Ⱥ=D=�.�=�ԍ=`��=ύ=P   P   �͜=㥎=/D=6Dʻ~��Hū�m�.��ԍ�4X���G��^����`.�$d��F<���4û&�D=���=�ڜ=���=���=P   P   |�=���=�~�=.D=� �vQ��[@v��ܾ����d0�µ���ܾ��u��뿽k�ۺXxD=ޤ�=6�=N��=&x�=P   P   �p�="��=���=⥎=��C=��<��a���Ych�@���
��,Uh���ĥa���<�7D=Qڎ=M(�=2Ǭ=_{�=P   P   ���=��=^�=�ǔ=��=1G:=PA�<�@M��C��񚽛-�����W�B���L����<B�:=}$�=�=��=
+�=P   P   	+�=t�=Bm�=�N�=t=�=��j=o�-=V �<af;�l���ͼ��ͼ��k�(j;���<v.=(yk=�{�=_��=���=P   P   ��=��=J�=wM�=�}�=�hw=ɸG=W:=b �<ƛ�;�ч� q���.�����;�<-�=�mH=�x=ƍ=_��=P   P   }�=nF�=H:�=�ǔ=�;�=fw=GL=�}=�ط<��<�t�V6����{���}�<�k�<uT=��L=�x=�{�=P   P   z$�=3��=NK�=�=<�=V�j=�G=Bz=��<��;,���,l������j�����#�;�Ҹ<tT=�mH=$yk=P   P   9�:=xP9=��4=��4=�_9={:=�#.=�F=4ҷ<�K�;B�������C|ԼU Լ>���q��#�;�k�<*�=v.=P   P   ܧ�<�n3< 2�:h*�\��:�6<���<A��<)X�<��<����Ꞽ
p�/����<�������}�<�<���<P   P   �L���'�畽�`½�½�����%��=G�{�s;O�;�a��l���Լ�?�.�P Լغj�Z���s��;b'j;P   P   q�B��)ܽ~�=�ꫂ�y.���I��ն<��)ڽ�g@�h9g��������VU����Լp�;|Լ��������.��+�k�P   P   ���	�2�&��������������_���t�0�"��.�ʼ�[������l�Ꞽ����l�E6�q���ͼP   P   �-���_����M_E�#E�����@㊿�VD�{�[]�5(��)�ʼ����oa�i����������1t��ч���ͼP   P   ���_�[���kx�d]ȿn� �r ��ǿ�v�����Y]�{"��M9g�~�;��<L�;��;�<国;�l�P   P   �C�R�2����*}x��"㿅M&��=���%�p��v�w�n�0��g@��s;7X�<Aҷ<��<�ط<m �<hf;P   P   �@M��*ܽ������E��ȿ�i&�S�W�J�W���%���ǿ�VD�X����)ڽx=G�T��<�F=Iz=�}=]:=\ �<P   P   RA�<y(�Y�=�Yn������1� �n=�P�W��=�m �:㊿���ɶ<���%�ڙ�<�#.=�G=ML=ϸG=s�-=P   P   4G:=��2<����䂾�!���/� ��i&��M&�i� ��������I�����46<{:=]�j="fw=�hw=��j=P   P   ��=&)9=���:��½P����!������ȿ�"�Z]ȿE����n.���½M��:�_9=D�=�;�=�}�=v=�=P   P   �ǔ=R�=F�4=T1���½�䂾Sn����E�}x�kx�@_E����߫���`½�*���4=�=�ǔ=xM�=�N�=P   P   _�=�3�=�?�=F�4=̫�:���S�=�~������L���������l�=��敽L5�:�4=RK�=J:�=K�=Cm�=P   P   ��=��=�3�=Q�=%)9=��2<r(��*ܽI�2��_�v_���2�u)ܽ��'��n3<�P9=6��=pF�=��=u�=P   P   ;ϒ=[]�=�a�=�ҁ=f(]=�=(&�<=!6��T$�.���h����̀��}$�ͬ6��<�=L>]=���=�o�=�d�=P   P   �d�=�]�=sp�=�͇=rx=j�R=A�=�|�<�ڻ;�>�(������8��I�;F��<=3>S=^Qx=�=˂�=P   P   �o�=5ύ=�^�=lɇ=ӏ~=��c=��>=R!=��<��E<*��;j.�:��;�F<���<��=�3?=K<d=W�~=�=P   P   ���=�W�=P�=ȁ=��w=��c=`�E=�=��<�ו<N%<�7�;2��;�&<k��<���<sL =�F=J<d=\Qx=P   P   F>]=�`=�0a=.�`=�]=��R=�>=�=���<��<@'$<ԯq;Z��:�uu;B�%<�=�<�3�<rL =�3?=/>S=P   P   ތ=�=G�=�=A/=�=]�=	 =�x�<��<�<S�:gJ���G����:L <�=�<���<��=�=P   P   e�<���;"�$�٧ʻ>?�<�;\�<���<"�<�ŕ<��#<C��:�������꠻���:C�%<i��<���<6��<P   P   �6��r����������m��2災����-2���;��F<m�$<��n;`M�c����G��uu;�&<�F<�I�;P   P   	~$�[�����P�D	f�+P�����趽5�"�-i����;"x�;B��:QM�����?J����:8��;��;�8�P   P   �̀��F�@Ɓ��H��<�辭��������q*���~�Ů��_z�:+x�;�n;���:��:�q;�7�;).�:���P   P   t��� 3�㮾�(���C�n�Y��C�����ح�:�1��(���������;y�$<��#<!�<Q'$<[%<(��;8��P   P   7���-�2�����+0��{��y>�����h���Q/��濾8�1���~�i���F<�ŕ<��< �<�ו<��E<�>�P   P   �T$��7��⮾�10��4���Qݿ%���ܿ礘��Q/��ح�m*�*�"�]��;"�<�x�<���<��<��<�ڻ;P   P   N!6��7���ā��6�0���jlݿ�M�>.��ܿe��������趽�-2����< =�=!�=V!=�|�<P   P   '&�<r4�̙��e����C��z���n���M�������C����������t�<d�=�>=d�E=��>=C�=P   P   �=���;���ɴP��A��HZ��z��flݿ�Qݿr>��d�Y����P�#災��;�=��R=��c=��c=m�R=P   P   h(]=�0=�G"�lզ�Fxf��A龪�C�-����4���{����C�.��3	f��m���=�L/=�]=��w=֏~=ux=P   P   �ҁ=��`=��=- ˻kզ�ƴP��e���6��10��+0��(��H���P�����#�ʻ%�=6�`=ȁ=nɇ=�͇=P   P   �a�= X�=xHa=��=yG"����ș��ā��⮾{��㮾7Ɓ�q��������$�T�=�0a=P�=�^�=sp�=P   P   []�=�͍=X�=��`=�0=���;k4��7���7�#�2��3��F��Z���r�M��;�=�`=�W�=6ύ=�]�=P   P   K�o=ݠl=<Fb=�M=�h'=VV�<~��;-ř�o�5��e���Ⓗ���8�5�|���P�;/��<zM'=~�L=)Eb= �l=P   P   ��l=l�l=�~g=�[= rF=��$=���<x�m<�XE�մe��벼����%f��L��Nm<Ј�<��$={�F=g�[=ȍg=P   P   'Eb=�,d=r4b=��[=��N=ʉ9=�I=�p�<���<��<�
;�k���;E=<q�<��<;|=��9=	�N=f�[=P   P   {�L=�WO=�OO=l�L=�YF=~9=��$=�*	=���<��<��8<s��;Tj�;_9<雑<6A�<i}	=G=%=��9=y�F=P   P   tM'=�?&=?W%=�:&=�='=h�$=79=�#	=��<��<��c<FB<�&�;��<Ee<r�<u��<h}	=9|=��$=P   P   ��<�a�<�ר<��<���<%�<:z�<�^�<���<ᣦ<U@j<��<��;�H�;��<Żk<r�<3A�<��<Ĉ�<P   P   EP�;~���V�b�+����La��ѕ����;{n<���<��<>�c<)�<<��;�+;a�;��<De<囑<h�<`Nm<P   P   0|���q1���������ݪ�yx��690�Ɉ��'+�ǟ<W�8<�<w�;��};�+;�H�;��<�^9<1=<��L�P   P   M�5�,f��Q����?���Q�Ba?�`N�G���^4���b��[;&��;��;w�;F��;��;�&�;Mj�;7�;&f�P   P   ������Vj�%���Ed˾2˾�����h��(��w��H������.��;"�<1�<��<MB<t��;�l����P   P   㒽��%������(����(���;�)O(��L��>왾B�$�5̑�D���[;a�8<I�c<`@j<��c<��8<�
;�벼P   P   �e��iv%��ҩ���M@n�^虿�Ù���m�w����@�$��w����b�ן<��<裦<��<��<��<�e�P   P   z�5�l��A���l��)���N̿Z�￬�˿Dņ�w�;왾�(��^4�]%+����<���<$��<���<���<CYE�P   P   8ř�~��X�i�����Cn�VX̿���S����˿��m��L��}�h�
G�������n<�^�<�#	=�*	=�p�<w�m<P   P   q��;��0����m~��Z�(�����&����S���Ù�#O(����XN�$90����;Gz�<;9=��$=�I=���<P   P   WV�<3y��Q����?��y˾ 	<����QX̿�N̿W虿��;��1˾6a?�lx��ѕ�%�<n�$=~9=͉9=��$=P   P   �h'=���<��`�}몽(	R��y˾W�(�|Cn��)��@@n���(�9d˾��Q��ݪ�pLa� �<�='=�YF=��N=rF=P   P   �M=zr&=o��<L��|몽�?�j~�����f�x��(�������?���������<�:&=p�L=��[=�[=P   P   =Fb=.vO=�%=o��<��`�N������P�i�:����ҩ�����Ej�E��v����b��ר<FW%=�OO=t4b=�~g=P   P   ޠl=<d=.vO=yr&=���<"y����0�w��e��`v%���%���f���q1������a�<�?&=�WO=�,d=m�l=P   P   ��/=*�,=^[!=�'=��<�`*<������j��W�������}��2�j�V~������(< ��< =�D!=�w,=P   P   �w,=Dx,=�'=@B=P�=?��<��l<j�:8yY�-VҼ �Y+���Ҽ5�Z�}X~:�)l<z�<F�=�;=ː'=P   P   �D!=��"=*A!=3=��=K��<���<�Ɉ<��;͒`�:�廡��滔�c�&�;���<3��<M��<2�=�;=P   P    =+�=m�= �
=x�=Ŗ�<���<p��<�a�<D�'<3��;�;GQ;p�;X6(<	��<չ<�*�<K��<D�=P   P   ���<K�<��<�Y�<��<�p�<�_�<3��<���<��i<��<��;��;�e�;s| <ܒj<C�<չ<-��<z�<P   P   ��(<�=�;ξG;��H;X��;U�)<c�l<~��<�R�<�i<�3<���;��;_c�;�C�;+�3<ڒj<��<���<y)l<P   P   �������A����]����<���r���؈:���;{�'<ѵ<���;���;�U�;��;�C�;o| <N6(<�%�;EV~:P   P   g~�-m�`c����ǽ�zǽp駽�_l�9�� 9X��wV����;�0�;EH�;�ܥ;�U�;_c�;�e�;[�;d�a�Z�P   P   H�j���н+�� :I�/�Z��H��H�˃Ͻwi�Ѽ
y��y;ں�;HH�;���;��;}��;$Q;B滩�ҼP   P   �}��5��uq�d���Ͼ$�ξ�J����p��}�t����?�����y;�0�;���;���;��;��;���e+�P   P   ����R\.�a�������0�#H�[i0�/���u���ǆ-�����?��x㻽��;ص<�3<��<0��;X���P   P   �W��K.�R���rA��􂿫��Uڰ�-���_������Ɔ-�q����ѼwV���'<#�i<�i<F�'<P�`�;VҼP   P   (j��	�Z���z7�SM���;��� �/� ��ᖿ]��r����}�mi��8X����;�R�<���<�a�<��;IyY�P   P   ����нm.q�gb���낿=�jOK�	*K�-� �*���'�����p�Ͻ.���و:���<:��<t��<�Ɉ<3�:P   P   �����l����펫���0�u���� �fOK��� �Nڰ�Ti0��J���H��_l�J��|�l<�_�<���<Æ�<��l<P   P   �`*<�h��$���H�� Ͼ�4H�s��
=�{;����t#H��ξ��H�d駽!���u�)<�p�<˖�<O��<A��<P   P   ��<'�;�`���Lǽh�Z�� Ͼ��0��낿KM�����0� Ͼ!�Z��zǽ������;���<|�=��=R�=P   P   �'=2��<��O;H���Lǽ��H�鎫�^b��r7�iA�֋��Y���:I�r�ǽ�]�U�H;�Y�<$�
=3=BB=P   P   _[!=<�=�1�<��O;�`��!򧽅��e.q�T���H���W����uq� ��Qc�������G;��<q�=,A!=�'=P   P   *�,=��"=;�=2��<-�;�h����l��н�	��J.�G\.��4��нm������=�;+K�</�=��"=Ex,=P   P   ���<���<&ֵ<j7�<��;c��ڼHmL�ދ��>껽M7ʽY���ז�XM��ۼUR��<�;Ծ�<���<_��<P   P   ]��<���<B��<j�<���<#�<�s��u����]�&�EyC���C���&��k�rKw�_�
�W�
<�L�<W߬<��<P   P   ���<�<ٖ�<-��<D��<�u<<
A�:�[ѻҬh�F����ɳ��ꢼFi�Z�һ�X�:I|<[su<�q�<T߬<P   P   ;�<�[�<1`�<!҆<Ad�<�u<M<�<��t;�c���ý�c����ཻﻺT�t;��<�L<Vsu<�L�<P   P   �<�;L��;F�;e��;l�;vO<�<��<�f�;�8m;���9���Ge6�y�����:fEn;���;��<=|<E�
<P   P   �R�N�
��Fހ��0M�7��5�r��:ܷt;M+m;jM;�=:+E�TW���:5�;WEn;-�t;�W�:Ξ
�P   P   -�ۼ-n!�cJ�<�Y���I�x� �˦ڼӨu���л�����<�9��
:q�'��P��V�շ��:N�:wﻺ��һ�Kw�P   P   jM�p���.ͽ��콷W�˷̽�����L�� 뼼�g�<+��y3���l�k����P��qW������ཻ#Fi��k�P   P   �ז��x..�˵Z��ul��`Z��-�)��"��"&�h�����,�6��l���'�7E�[e6����ꢼ��&�P   P   e����#��L���[���ھ��پ񴾙܀�&#��;����B��������a3����
:�=:���n��ɳ���C�P   P   X7ʽ��>�+������J8=�vW��<��+� 	����=�D[ɽ��B�d��/+��p=�9wM;���9Ľ�Q���QyC�P   P   G껽��>����J'����R�ȿuZȿa���Ҳ&�zn����=��;��&���g�G���f+m;�8m;�c���h�f�&�P   P   勖��#�B����<'�.�����H�B��L�$.��в&�	��&#��"��� �w�л�t;g�;��t;�[ѻ���P   P   OmL���!���v�Z�������{���z��L�]����+��܀��(�L���u����:��<�<�@�:�u�P   P   ʎڼ������-��$���=���ȿ/�B��{�?�B�jZȿ�<�����-�w�����ڼ�5��<M<<�s�P   P   n��	� ���̽T`Z���پ�}W��ȿ�����D�ȿ�uW���پ�`Z���̽j� ��6�O<��u<�u<#�<P   P   ��;йK��BI�J
��@l���پ�=�T���$������=8=��ھ�ul��W콊�I�h0M���;Hd�<H��<���<P   P   k7�<C�;.��O�X�I
�Q`Z��$���v��<'�
J'�����[����Z���(�Y�/ހ����;)҆<1��<l�<P   P   'ֵ<7�<Ӎ�;,���BI���̽��-�!��;������!����L��l..��.ͽOJ��	��UF�;9`�<ݖ�<D��<P   P   ���<�L�<7�<C�;˹K�� �������۟#���>���>���#��c��n!��N����;�[�<�<���<P   P   
<�K�;���;p��¸/�4|˼��2�@M��ɐ��f0ٽ���xaٽ�ൽW����3�j�̼�]1�ʦ��R��;`��;P   P   [��;���;�]�;	Ht;�����Қ��[ ��'6�ؙd������#�d�#�6�1� �d���3l���4�q;���;P   P   C��;��;p�;�>s;@c�:j���0�껠�d�T���Ğ�f0��P����5����e��컅�����:"�q;P   P   =����o�������"��NR���Xt�[�ݻ��0�ILw�rޙ�Y��Lj�����n�w�H(1���޻��v�����c��P   P   ^1��N��Y��M���0�ݲ��?�{�ݻ['��B���x=�'Y���c�]-Y�7�=����1���
�޻��Fl�P   P   }�̼8����M
��5
�� ��]�˼���y�d�`�0�M�����-w%�Iw.�o.�Ff%������S(1�Ěe�s���P   P   �3�kh�T��'���G'����g���2��P �����ew��_=��p%�L�����9�Hf%�?�=�}�w��5��;� �P   P   `��������i�P�n9���뽠��a*��v�5� 3�g�����X��q.������o.�e-Y�����/�6�P   P   �ൽ���;9:��vd��;u�1'd�L�9�Vb��.���d���
�� ��&�c��q.�L�Lw.���c�Tj��	P�1�d�P   P   �aٽ��/��愾Hĵ��
ؾ��׾/a��T~��EJ/�ǌؽh&���� ����X��p%�.w%�'Y�$Y������P   P   ��}HI�+ꧾ���x5��M��%5��[�X����H����g&���
�d����_=�����x=�wޙ�l0���P   P   p0ٽ�4I�U���p!�܆�<��0	��烆��� �v�����H�Čؽ�d�3�]w�I��B��PLw�͞��d�P   P   А���/�j̧�kd!�߮��'�
���.���
�E<���� �X��BJ/��.��q�5�����W�0�U'����0�Y����'6�P   P   EM��N���������cІ�w�
�nQ_��#_���
�テ��[�P~��Rb�\*���P �l�d�m�ݻX�ݻ��d��[ �P   P   ��2�,����9�;���R\5�C����.�iQ_���.�'	���%5�'a��D�9������2�����?��Xt�0�껊Қ�P   P   7|˼Eg�2��5d���׾:�M��B��q�
��
�<��ރM���׾&'d����u�g�N�˼̲�R��P����P   P   ĸ/�\>��懽���u���׾N\5�^І�֮��܆�x5��
ؾ�;u�f9�>'��� ���0�g"��pc�:���P   P   p��gJL�w�	�A�����2d�7������cd!��p!����=ĵ��vd�P�����5
��M�j���>s;Ht;P   P   ���;~ߨ�AXW�v�	�~懽/����9�����ç�U��"ꧾ�愾/9:��i�
T��~M
�lY�n�����;�]�;P   P   �K�;	��;ߨ�fJL�Y>��Eg�,��J���/��4I�rHI���/��������Zh�!����N�}o��'��;��;P   P   a������F�lg����߼C''���o�7��?6̽qV� ��� �콪�̽�h��
+p��'���༻��g�G�V��P   P   Y��w���f(�ۺV����$�ͼ�P���=��yo�5����������;0��}�o�AI>����`SμyU��K�W�|�(�P   P   n�G�Q�B�o=G��V�|w�������� ��2��;8/�ϋB���I�F�B�jx/�O���G񼚔��6����w�O�W�P   P   ���Dn��sX���Γ�����b����ס��ɵ�5�м�W����>�9J������
CѼ�<���J��9��~U��P   P   ���)�１2��
f�.p�X�ͼ����е�7���������ɼQӼ��ּ�eӼ�ʼzվ��ⶼ�<������jSμP   P   ��'���=��K�R�J�O�=�\'�eg�F����м����G��`t��΅��:�������
n��|վ�CѼ�G���P   P   +p�H'��{.��J��T��������o�{�=����1���ɼ�k��N�������$�������ʼ��V��KI>�P   P   i��ݹҽ�����F�}����6ҽ���1o���.����=%Ӽ6t���������<����eӼ���rx/���o�P   P   ��̽��"�;�E`���n�� `��?;�����˽����:,B��H�ּ6t��O��Ѕ����ּ=J�O�B�B0��P   P   �콽m2� �� è�͋ľ5iľ{q��W�S�1����<���/I��<%Ӽ�k��bt��QӼ�>���I�����P   P   ���тH��S��Ss�~��a�*��Y���羧ڜ���G�K���<��9,B������ɼG����ɼ��֋B�����P   P   {V�qH��3��h]���X�AV��7���ZX���
�9�����G����������.��1��������W�@8/�:��P   P   F6̽-?2��:��tT���v��¿��� ����v���
��ڜ�P�1��˽�1o�����м6���8�м5���yo�P   P   <��3��v���I農�X��¿�T��9������ZX����	W�����v�=�?��е��ɵ����=�P   P   ��o��Bҽ�[;�[���t���[��|���T���� 7���Y�uq���?;��6ҽ��o�`g�����ס������P�P   P   E''��������!�_��jľ"�*��[��{¿�¿9V��W�*�,iľ� `�r��������['�P�ͼ^������%�ͼP   P   ��߼�J=�+ƣ�~��nn��jľq����X���v���X�u��ľ��n�?�L��F�=�$p༮���ww����P   P   lg�����V|J�G諾}���_�W���|I�nT�`]�Fs�è��D`����I��G�J��e＝Γ� �V�غV�P   P   ��F��Δ�kY��U|J�)ƣ�|����[;�o���:��{3���S�����;�y��q.���K��2��kX��f=G��f(�P   P   ��'(B��Δ�����J=������Bҽ/��'?2��pH�ǂH��m2���ѹҽ@'����=���<n��I�B�s��P   P   ���0�ɼ@��|����,��-_�� ��)���^ٽߚ��l������4�ٽ�k���N����_�a-�q��Q���ɼP   P   ��ɼ�ɼ�Լ
���0�R�#�ÝG�!3r�����������0����ݡ�9J��U�r��H���#�;��'C뼔aԼP   P   Q�k��'%�m���&��^�	��[���1���J�6.b�es�F@y��,s�Npb��(K��B2�ү�K�	�W���*C�P   P   t��@�	�T�	�����L�ː	�@����!��A-�^�7��=��=�V�7�zw-�K^!�\S��>�M�	�=��P   P   g-�34�۰6�d�3���,�ϰ#�g������'�������q����Q��JV�f��]S�֯���#�P   P   �_��At��#�������s��Z_��G���1�7!�I!��A�_��`)��/�����c�KV�N^!��B2��H�P   P   �N��2ɦ��������g��������T"r�]�J�+-�q������al�����S��~w-��(K�^�r�P   P   �k���v߽������s���b��߽!����[�a�ݎ7��p����e�al��/���[�7�Vpb�?J��P   P   >�ٽdg�3�3�d�P��6\�+�P��3� ��ٽ
u��5�r�<�=�o������a)�s���=��,s��ݡ�P   P    ���mU,�0�i�������U����I���%i�,�+�
��`4����x�;�=��p����`������=�N@y�7���P   P   v���(>����Q����<�&��#��m������=�S:��`4��3�r�܎7�q��A����a�7�ls���P   P   ����>��ړ���߾Ȼ�$XB�a5B�Pu��i߾�}���=���u��X�a�+-�I!��'��A-�<.b����P   P   �^ٽ�.,������߾�`.��.w��Ō���v�*	.��i߾���)�+��ٽ�[�J�6!���!���J����P   P   -��M4�(ti���������2w�A/��D����v�Mu�|m���%i������O"r���1�������1�%3r�P   P   � ���߽%�3�Ld��*%�_B��،�?/���Ō�[5B����I����3��߽����G�g�@���[�ƝG�P   P   �-_��m���V���P���������_B��2w��.w�XB� ��N���#�P��b�����Z_�̰#�ʐ	�]�	�S�#�P   P   ��,���s��1����\�����'%򾧳��`.�����<�����6\�m���f����s���,��L��&���0�P   P   |����3�����q������P�Id��������߾u�߾G������Z�P����������^�3����j��	��P   P   @�⼁J	��K6�����1���V�"�3�"ti�����ړ����$�i�)�3���������#��հ6�P�	�#%��ԼP   P   /�ɼ>t༁J	���3���s��m���߽J4��.,��>�>�dU,�]g��v߽*ɦ��At�-4�<�	�g���ɼP   P   �%�f��'*�?�?�Gm`�^���T��S[����޽>���[�������6߽����g���Æ���`�n@�5\*���P   P   �����6#�=.�r?��&X���w��Z�����K���ϑ��P�������[/��H���]x�ӈX��?��A.�&[#�P   P   7\*�	)�LE*�'.��95���@��MP���c�b:y�\���3���94��Ũ������I�y�9d���P�!�@�py5��A.�P   P   q@���@�a�@�;�?��?��@��D���J�X�S�Qg]�[�e���j���j��f�֠]���S���J�JjD�"�@��?�P   P   ��`��$g��wi�3g��`�=?X��UP�K�J�&H��"H�h�I���K�|tL��K�a�I��YH��FH���J���P�׈X�P   P   Æ��Ï�!���j锽����U���|�w�N�c���S�H��"A��=��
<��<��=��NA��YH���S�9d�#]x�P   P   m���6���ݰý�Ƚ��ýz��iV���Q���y�nN]���I�g|=��6�j�4�O�6��=�c�I�ڠ]�O�y�L���P   P   ����=��6�.#
�~
�������@���ޠ�Cd����e��K��;�&�4�j�4��<��K��f����a/��P   P   �6߽�C��P'���<��5E�n�<��'���
���޽�Z��.j��˝j�|JL��;��6��
<�tL���j�ɨ������P   P   ������!�H�N��"z�P���������y���N��3!��t��wA������˝j��K�g|=��=���K���j�=4��V���P   P   d��Y�.�vn��%��̹��&ƾ+����㚾��m��.�ɂ��vA��.j����e���I��"A�j�I�_�e�7���ԑ��P   P   E����.�0�z�ײ��a�㾡Q�A��c㾍a��z��.��t���Z��Bd��mN]�H��"H�Tg]�_���P���P   P   ��޽�o!�\n���������a�b7+��?������a����m��3!���޽�ޠ��y���S�&H�Z�S�e:y����P   P   W[��0��N�\����xc�e)=�=��?��c��㚾��N���
��@���Q��L�c�J�J���J���c��Z��P   P   T��M��d '���y�ཹ�:U��G+�c)=�_7+�A�%�����y��'����eV��x�w��UP��D��MP���w�P   P   _����d��	���<�{����+ƾ9U�uc��a��Q��&ƾ�g�<����y��R���:?X��@���@��&X�P   P   Gm`���xcý��	��E�z���ݽ��z�㾈��X���˹�J����5E�y
���ý�����`��?��95�r?�P   P   ?�?���f�Ƿ���Ƚ��	���<���y�X������Ѳ���%���"z���<�)#
��Ƚe锽-g�8�?�&.�=.�P   P   �'*��W@��i�Ƿ��wcý	�b '��N��[n�&�z��un�?�N��P'��6�հý���~wi�]�@�JE*��6#�P   P   f���(��W@���f������d��I��-��o!��.�R�.���!��C��=�/����Ï��$g���@�)���P   P   �L���O�{[���n�P���y���2���ȯȽ��߽��'	��4���$���Ƚ��E䘽W҅���n�N2[���O�P   P   ��O���O�Q�T���^��Yn���� ���q���E��kӺ�s����½��cp��4���Տ�o6����n���^��T�P   P   O2[��Z�[�-�^�p?e�Jo�2�|�K̆�S���~֗�����ʽ��'���a�ڏ�����~N}�ԗo��e���^�P   P   ��n�7Bo�55o�h�n��ln��Po��Ar�Άw�ث~�b@������ř�����������\����~���w�r�՗o���n�P   P   Y҅���������v������s����|�f�w��it��s��3t��5u���u��Ku��\t�)�s�رt���w��N}�q6��P   P   I䘽%p��)��������S��S���{����Ɇ�E�~�!�s�QGl��h�4Nf�'Xf��9h��xl�*�s���~������Տ�P   P   ��<���1�ʽ��νs�ʽ�Q��3���A���8����3��� t��h�Va��5_�ja��9h��\t��\��ڏ�4��P   P   ��Ƚ�=余r���u��k��:�����v�ȽR*������֋��Eu�4:f��,_��5_�)Xf��Ku�����d�gp��P   P   �$�H����a})�JC/��`)����?�߽¢���v��!{��x�u�4:f�Va�5Nf���u� ���*�����P   P   <��0��L6�/PS��e��e��S���5�
��X~��������!{��Eu��h��h��5u�Ǚ��ν���½P   P   .	���n�ȋK��z�����n떾���w�y�X7K��(�w�������v��Ջ��� t�QGl��3t���������x���P   P   ��f��S�u��O���Om��B\��<y���݈�gRS��(�W~����������3��!�s��s�c@���֗�oӺ�P   P   ��߽���zK��	��L���Ӿm�ᾐkӾ��݈�V7K���=�߽Q*��7���D�~��it�ګ~�U����E��P   P   ˯Ƚ2)���5� �y�����Ӿ�8�*�kӾ:y��t�y���5��s�Ƚ?����Ɇ�f�w�φw�L̆�s��P   P   4�����㽏��R0S�ϥ���p���ᾡ8�i��>\������S������1���y�����|��Ar�2�|����P   P   z����A���+��\)��e��햾�p���Ӿ�ӾJm��j떾�e��`)��:���Q��Q���q���Po�Jo����P   P   P���d8��Stʽ>W��-/��e�Υ�����G��J��������e�DC/��k�n�ʽ�S�������ln�o?e��Yn�P   P   ��n�gY������&�ν>W� \)�P0S���y��	��q���z�'PS�[})��u���ν�����v��f�n�,�^���^�P   P   {[�$o��Z������Rtʽ�+�������5�zK�ڦS���K�E6�����r��+�ʽ%������25o�[�P�T�P   P   ��O�*�Y�$o�fY��c8���A�����0)�����f��n�+��H��=�6���!p������4Bo��Z���O�P   P   -�v�r�y���������hۖ�ӯ��C����̽h�޽�G�V��8[���޽�ͽIt��rަ����+��������y�P   P   ��y��y�rE~�w��������ԓ�~1������跽����yQǽ�ZǽO������㫽�\��m�����5���g~�P   P   ������p���������/����ѫ����v������9ɫ�l)��,�������җ�D落�������6���P   P   -���dՊ�"ϊ�n���񋊽��&"��C������4���ܖ�h���m����O���>���g��G������P   P   ���H?�����1���ꖽ�ۓ�\��A��׬��������?��Fb���I�����_!��=Ќ��g��F落o���P   P   uަ�r ���w���n��謽g����2��z���l����ށ��gg���s���x��?v������`!���>���җ��\��P   P   Mt����Ž�yν�ѽ�bν��Ž�B��Q���Z瞽+(��Z���9b���.��(���8��?v������O������㫽P   P   �ͽ�+b��L���=���7�,��{�̽.ѷ�
i��dȖ��/��Ti��!#��(���x���I���/������P   P   ��޽,z���'�����������*���z޽י��c����K���L��Ti���.���s��Gb���m��o)��S���P   P   >[���}�!��45�Ѻ@�G�@�5��}!�<�
��	뽓ǽ	����K���/��9b��hg��?�� h��<ɫ��ZǽP   P   [������0��N���d�"xm��d�d�M���/�����ｓǽb���dȖ�Z���߁������ܖ����}QǽP   P   �G뽱���l5���\�o��z���p��NW��Ѣ\��55����	�֙��	i��+(��������4��x�������P   P   l�޽J��	0�'�\��ȅ�(]��:���rL������Т\���/�;�
��z޽,ѷ�Y瞽l��׬��������跽P   P   ��̽�K���!� �M��k���]���i���b��rL��MW��b�M��}!��*��y�̽O���y����A��C��ҫ�����P   P   C��r��\�#5�!�d��{��G����i��8����p���d� 5���(���B���2��[�&"������1��P   P   ԯ����Ž�,�/��^�@��ym��{���]��&]��	z��xm�C�@�����7󽳝Že����ۓ���.�ԓ�P   P   iۖ��Ҭ��GνC��	��^�@��d��k���ȅ�o����d�̺@����=���bν謽�ꖽ�����������P   P   ��������M��rѽC��.��"5��M�#�\���\��N��45����L���ѽ�n��|1��l�������w���P   P   ��������w왽�M���Gν�,�[��!��	0��l5��0�y�!��'�$b�yν�w�����!ϊ�o��qE~�P   P   r�y�s����������Ҭ���Žo�ὲK��H���������%z��	���Žo ��F?��bՊ���� �y�P   P   ����Lm��Eƒ�����]���>�������Ͻ�rܽ���b2齗��*�ܽ�1Ͻ���e��뀤��4���ْ�>w��P   P   >w���r��Y���7��H��㡽u1���8��Ǿ� aƽu�ʽ��ʽ
uƽ�侽�\���V������7��;O��Nh��P   P   �ْ� ]���Β��;������y���P�������Ӫ�������������;����X��t�������ݖ�<O��P   P   �4��H��mB��%�����{���v��-'��Re��Zϡ��ߣ����&���衽����I�����������7��P   P   퀤�cI���즽=��\i��(衽?Q���%��k���P�G����Κ�����ٚ�GӚ�g���Λ�I��t�����P   P   �e��TE����������0���F��>1��N���`���횽ė��˕��ߔ��䔽8ڕ�2ۗ�h������Y���V��P   P   
��Q�ɽPнN�ҽ�=н��ɽ���0��Ȫ��á�u����ƕ��䒽����V9ڕ�HӚ�衽�񪽍\��P   P   �1ϽY߽�����	󽽿���޽��ν�����ﯽ}ͣ�V����Ք��������䔽ٚ��=���侽P   P   /�ܽ���0��.������������BTܽ�@ƽ����@����̚��Ք��䒽�ߔ�����(������uƽP   P   ���:t���Y,��&��&���U��R����	tʽɴ�@���V����ƕ��˕��Κ�������ʽP   P   g2齫A���!6/�:w=�J�B�d=��/���������tʽ����}ͣ�u���ė�H����ߣ�����x�ʽP   P   ���-=��N�\�8��UN��5[�+[�:N�)b8�Y*�����彫@ƽ�ﯽ�á��횽P�[ϡ����#aƽP   P   �rܽ>h����Ԃ8��T���i�V�q���i�=�T�)b8����R�ATܽ����Ȫ�`��k���Se���Ӫ�Ǿ�P   P   �Ͻ����
��+/��QN�`�i�8=z��5z���i�:N��/�S�������ν�0��N����%��-'�������8��P   P   ������޽������o=��6[���q�7=z�T�q�+[�d=��������޽��<1��>Q���v���P��v1��P   P    ?��Q�ɽ���1��&�l�B��6[�^�i���i��5[�G�B��&�����뽪�ɽ�F��'衽{��y��㡽P   P   �]��* ��L)нL��-���&��o=��QN��T��UN�6w=��&�����	��=н�0��Zi���������H��P   P   ���K*��j۸�ٍҽL��0����+/�т8�X�8�6/�V,�.���J�ҽ ���=��%���;���7��P   P   Eƒ��0���Ҧ�j۸�K)н�������
����}N�����-�����Pн~����즽lB���Β�Y��P   P   Lm���N���0��J*��* ��P�ɽ��޽���<h�+=��A�7t����U߽M�ɽQE��aI��H��]���r��P   P   �|�������W��Oi��DƮ������Ľ�н[ڽ��Ru��&,ڽB,н�Ľ�/���⮽À��Eh��6���P   P   6������jR��۔��w���Ь��F��M+��?�ý�bɽa�̽۟̽�rɽ��ý
I���e��﬽����R����_��P   P   Eh������^������ả��Φ������E���⳽�m��������ú���1���Qc��Mު�w립ӣ�S���P   P   Ā������ɂ���r��_{��#Ц�$���������o�����������w)�����ͪ�������x립����P   P   �⮽�F���ư��;���ή�lԬ�e���l򨽄�����ԧ��̛��ϟ��Ϥ�����
��6ȧ����Nު�	﬽P   P   �/��h���I������鼽���F��!B������:-��gn��c���Ş���{���A��
��ͪ�Rc���e��P   P   �Ľ��˽ ѽ�ҽ��нu�˽&�Ľ$��;س�����ɟ��0j��퟽d�������{��������3���I��P   P   E,н�
ܽ�t�U�꽖��I\�f�۽�н��ý�ݷ����Ď��r������d��ƞ��Ф��x)������ýP   P   ),ڽ N�~��t���m����Z��v!뽔�ٽ�Hɽ!����쮽ҍ��r���퟽d���П������ú��rɽP   P   �Pp��%���t�q�k��d�����>����ེw̽�����쮽Ď��0j��hn��͛��������ޟ̽P   P   Uu�y1���-����#�rl&��#�����������I㽺w̽!������ɟ��;-��ԧ�����o���c�̽P   P   ��<+��@��F����-��t5�Kn5�ʏ-�Z���q���������Hɽ�ݷ��������p�����bɽP   P   ]ڽ�^���'����w1��>���B��>�e1�Z�����>����ٽ��ý:س�������������⳽A�ýP   P   �нb3뽡�������-��>�Z�G�u�G��>�ɏ-�������t!��н$�� B��l򨽓󨽧E��N+��P   P   ��Ľ��۽gb���j��#��t5�9�B�Z�G���B�In5��#��d��Z��d�۽$�ĽF��d���$��������F��P   P   �����˽�V�`}��i�2l&��t5��>��>��t5�pl&�k���F\�s�˽���kԬ�"Ц��Φ��Ь�P   P   DƮ�]ݼ���нS��~e��i��#��-�w1���-�#��p��m���꽵�н�鼽�ή�^{��ả�w��P   P   Oi��-��l����ҽS��`}��j�������D������t�q��Q���ҽ����;���r������۔��P   P   �W��Zt��:���k�����н�V�eb������'�>���-�"��~���t� ѽG���ư�Ȃ���^��jR��P   P   ����*�Zt��-��\ݼ���˽��۽`3뽨^��8+��u1��Lp���M뽰
ܽ��˽f����F������������P   P   Z-��|*��x'�����鿶�Ҿ��ǽ�_н��׽��ܽ2�޽B�ܽ)�׽�uн��ǽ�뾽�ֶ�&��=5���1��P   P   �1���-�����?2���(��o=�����;����ƽ�I˽>�ͽ��ͽ_V˽��ƽT���5���V��S?���C�����P   P   >5��S٪�v-���4��*����y��ޞ��)-���º��ݽ�������������׺�F������ᑰ�����C��P   P   &�� "��������,��z���"��+-��S����紽��������Ŷ�z ������홳�G���<��ᑰ�S?��P   P   �ֶ�g淽�E��Oݷ�8ƶ�@��Z���I,������o��T�����T������.�����u1�� G�������V��P   P   쾽���=kýfýD����վ����)���}��3m���!������I髽6�N����3�����홳�F���5��P   P   ��ǽ}Jͽe	ѽwZҽ*�н�5ͽ��ǽv5��ݹ��1ߴ�K�����������ة�����N����.�������׺�T��P   P   �uн�Iٽ�,�M��a����.ٽ�Uнf�ƽϽ��������᫽�ԩ��ة�6����{ ������ƽP   P   +�׽{q�9R�_���<e��1���8ｦO���׽ 5˽1鿽%����򯽝᫽����I髽U���Ŷ����aV˽P   P   D�ܽt'�y���K�N��N��t@��Y������ܽݘͽL���%����������������������	�����ͽP   P   5�޽���0���_��[�!���S��Q�y��B���޽ݘͽ1鿽��K���!��U��������@�ͽP   P   ��ܽ����[�Q� �~�i��� B�	K�A����ܽ5˽Ͻ�1ߴ�3m���o���紽�ݽ��I˽P   P   ��׽D���JO�	���t"��M%�Kn"���� B�x������׽f�ƽܹ���}�����T����º���ƽP   P   �_н=]�zj��	[�Q��t"��K(��I(�Jn"����Q��Y���O佭Uнu5���)��H,��+-��*-���;��P   P   �ǽ�1ٽI>�ID�@X�(�JP%��K(��M%�h��S�r@�8�.ٽ��ǽ
��Z����"��ߞ����P   P   Ҿ��1ͽ��԰��+����(��t"��t"�|� ��M��/����཯5ͽ�վ�@��z���y��p=��P   P   鿶����]�н���>Z��+��?X�P��� ��[�L��9e��^��(�нC���7ƶ�,��)����(��P   P   ����ѷ�Wý�Hҽ���Ӱ��ID�[�IO�Q��_��K�[���J��uZҽfýNݷ�����4��?2��P   P   x'��J���5��Wý\�н��H>�xj�����[�.���y��6R･,�b	ѽ;ký�E�����u-�����P   P   |*��YϪ�J���ѷ�����1ͽ�1ٽ;]�B�������q'�wq佂Iٽ{Jͽ���f淽�!��R٪��-��P   P   �{���G��{���ܖ���Լ�6ý�ɽ�Xн��ս*�ٽd�ڽ��ٽL�սjн
�ɽ�&ýe缽���������M��P   P   �M��J��,`������ޱ��9���I?��1�Ľ�7ɽ݃̽�Qν,Uν�̽�Gɽ�Ž�T��/ǻ��ķ�]���di��P   P   ����m��:��������������|s���4��}�|N½p�ý|ĽO�ý�[½����I����������]���P   P   �������o��������������>����Q��8T��"_��%=��$�������
G���n��Ch���g��K�������ķ�P   P   f缽鲽�m���e���ټ� ���s���P���p���޷������n��2j��*u�������𷽫����g�����/ǻ�P   P   �&ý7XŽ��ƽh�ƽLŽ�ýX>���1���P��Gܷ����������#��'���ȴ�C����Dh���I���T��P   P   �ɽ�ν�н(�ѽ�н#�ͽ��ɽ��Ľq쿽HX��ɉ������W���y��/���ȴ������n������ŽP   P   jн��ֽH�۽j�޽B�޽�۽b�ֽ�Pн%-ɽHB½�1��1e��
��v���y��'��*u��G���[½�GɽP   P   N�սZ߽��潻*�-�I �l�� ߽��սys̽��ý쭼��\��
��W���#��2j������P�ý�̽P   P   ��ٽ_�g5�X���\=���7��I���o��C彵�ٽ'<νgĽ쭼�1e�����������n��%���|Ľ.UνP   P   f�ڽ8����6)��/����*�K�i�����ڽ'<ν��ý�1��ɉ����������&=��q�ý�QνP   P   ,�ٽG��׼��C��#�	��������	����6����轵�ٽys̽HB½HX��Gܷ��޷�#_��}N½߃̽P   P   ��սU彍|������F�d�D6��_�-?����~i���C���ս%-ɽq쿽�P���p��9T��~��7ɽP   P   �Xн
߽;*��%��	��c���K��_��	�J�n� ߽�Pн��Ľ�1���P���Q���4��2�ĽP   P   �ɽh�ֽ@�潏���l-�8���7���D6�����*�H���j��a�ֽ��ɽW>��s��>���|s��I?��P   P   6ý.�ͽ=�۽��6�����8���c�d�������7��H ��۽"�ͽ�ý������������9���P   P   �Լ�;EŽ[�н��޽f��6��k-��	��F�"�	��/�Z=��+�@�޽�нLŽ~ټ��������ޱ��P   P   ܖ��9����yƽ׺ѽ��޽�콎����%����B��5)�V����*�g�޽&�ѽg�ƽd��������������P   P   {���L����뽽�yƽZ�н<�۽?��:*�|��Լ������e5����F�۽�н��ƽk���n���9���,`��P   P   �G���d��L���9���;EŽ-�ͽg�ֽ
߽U�E��6��_�X߽��ֽ�ν5XŽ貽����m��J��P   P   �Ϸ��q��vU��e��(u��Q<ƽtS˽�3н<HԽ�׽��׽Z׽aRԽ�Aнc˽�Lƽk����q���^���v��P   P   �v��t���Q��|�����������Ľ��ǽ=�ʽUͽ�ν��ν8]ͽ��ʽ\�ǽ,Ľ��������T���Y��P   P   �^��!��MY�����.��z������U�����ý�Ž>�ƽpCǽ��ƽ�Ž��ý[���{���Vн�o<��U��P   P   �q��Xf��=c��fi�����������,���˾�I����S������S���V��&����`�������ݾ�?��Vн�����P   P   l����½_L½t½�x����������˾�C������1Y���8���0��Y>��d�������*���ݾ�{�������P   P   �Lƽ@�ǽ��Ƚ\�Ƚ��ǽ�=ƽ�Ľt���B���}������$��k���(����'���+����������[���,ĽP   P   c˽$vνłн�8ѽ�{н�hν�Q˽�ǽ�ý	N���T�����'���gL���Ź��'��d���`����ý]�ǽP   P   �Aн�սD�ؽ�ڽ�ڽx�ؽ� ս�-н��ʽW�Ž�����0��ܚ���I��gL��)���Z>��'����Ž��ʽP   P   bRԽ�۽"���e�X���]佥�ག�ڽ-=ԽHͽ@�ƽmG��&��ܚ��'���k����0���V����ƽ:]ͽP   P   \׽�߽*H�2�Re�ja�{&��6�jx߽M�ֽ �ν2ǽmG���0�����$���8���S��qCǽ��νP   P   ��׽������%��s��gb��ik��$�󽶦���Ὢ�׽ �ν@�ƽ�����T�����2Y�����?�ƽ�νP   P   �׽���F�Y�������,��f��"��������5����M�ֽHͽV�Ž	N��}��������S���ŽUͽP   P   =HԽy�߽W�뽏���U� ��B��v��?�U� ��������jx߽-=Խ��ʽ�ýB���C��I�����ý>�ʽP   P   �3нC�ڽ�?�;������B�Ŷ�Ƶ��?�"���$���6罁�ڽ�-н�ǽt���˾��˾�U�����ǽP   P   uS˽�ս��^*�<o��
���w�Ķ��v�e��hk��z&���� ս�Q˽�Ľ�����,������ĽP   P   R<ƽ�fν}�ؽY\�>`�a��	���B��B�,��eb��ia��]�w�ؽ�hν�=ƽ��������z�������P   P   (u����ǽ�uн��ڽ-��>`�;o�����T� �����s��Pe�V���ڽ�{н��ǽ�x������.������P   P   e���½��Ƚ�.ѽ��ڽY\�]*�:�󽎗��W���#��2��e��ڽ�8ѽ[�Ƚs½ei�����|��P   P   vU��\���B½��Ƚ�uн|�ؽ�ཾ?�V���F���(H�!��C�ؽĂн��Ƚ^L½<c��MY���Q��P   P   �q�����\���½��ǽ�fν�սB�ڽx�߽�Ὑ���߽�۽�ս"vν?�ǽ�½Wf��!��t��P   P   b������	~������{�Ľ�ȽXh̽�н�	ӽlս��սrս�ӽн�t̽ѣȽ�Ž>��������	��P   P   �	���������
�������VĽ��ƽͫɽ�̽F�ͽi�ν��ν��ͽ̽B�ɽǽidĽ�½ ��U���P   P   ����$T�����Z��*����*½!�ýb>Ž�ƽO ȽoɽhVɽ�ɽ�(Ƚ	�ƽPLŽN�ýb8½3�����P   P   ?�������r���l���A���+½�½	�½N�ý�ĽƑĽB�Ľ��ĽV�Ľ3%Ľ��ý�ýT�½b8½�½P   P   �Ž�pŽ �Ž�kŽB�Ľ0WĽ��ýR�½�n½�½G���V���ŧ��,���)���<½<}½�ýN�ýidĽP   P   ңȽ+�ɽ_�ʽ�ʽ��ɽ;�Ƚ*�ƽ+<Ž�ý2
½g�����4���u������k���<½��ýQLŽǽP   P   �t̽��ν|>н�н�8нޱν�f̽�ɽ��ƽ�Ľ�������K���W���)�����)���4%Ľ
�ƽC�ɽP   P   	н؝ӽIֽ_�׽��׽�@ֽِӽ н{̽�Ƚ%�Ľ�������$���X���u���,���W�Ľ�(Ƚ̽P   P   �ӽ6�׽Uܽ�޽��߽��޽z�۽��׽Fӽ��ͽ(�Ƚ �ĽY�������K���4���Ƨ����Ľ�ɽ��ͽP   P   sս�=۽-��L�佗;��8������o.۽��Խ"�νIɽ �Ľ��������W���B�ĽhVɽ��νP   P   ��սzݽ���&��?��{���%�齯��^�ܽ�ս"�ν(�Ƚ%�Ľ����h���G���ǑĽpɽj�νP   P   mս8 ݽ�
�AG�+��Ͽ������ٿ�<�<��^�ܽ��Խ��ͽ�Ƚ�Ľ3
½�½�ĽP ȽG�ͽP   P   �	ӽQ8۽c��F콢A������������:�<콯��o.۽Eӽ{̽��ƽ�ý�n½N�ý�ƽ�̽P   P   �н��׽��ཌ��o������W>��{<�����ؿ�$���ཱུ�׽н�ɽ*<ŽQ�½	�½b>ŽͫɽP   P   Yh̽-�ӽ��۽���*����������V>���������������y�۽ؐӽ�f̽)�ƽ��ý�½!�ý��ƽP   P   �Ƚw�ν�?ֽޯ޽8罫��������������ο��z���8罷�޽�@ֽޱν;�Ƚ/WĽ+½�*½�VĽP   P   {�Ľ��ɽS4н��׽̡߽8�*��n��A�*��>��;罶�߽��׽�8н��ɽA�Ľ@���*�������P   P   ����tfŽyʽl�н��׽ޯ޽��佋��F�@G�$��K���޽^�׽�н�ʽ�kŽl���Z���
��P   P   	~�������ŽyʽS4н�?ֽ��۽���b�㽏
彯��,��SܽIֽ{>н^�ʽ�Žr���������P   P   ���[O������tfŽ��ɽw�ν-�ӽ��׽P8۽7 ݽxݽ�=۽5�׽֝ӽ��ν*�ɽ�pŽ����$T�����P   P   �����R½�sý�BŽ[�ǽ�Zʽ�4ͽt�ϽҽV�ӽ�Խh�ӽҽ_�Ͻ�>ͽ�dʽ��ǽKŽ9zý�U½P   P   �U½FT½��½@�ýOZŽ�*ǽ�*ɽ+˽��̽�Jν�Ͻ�Ͻ�Oν<�̽�4˽76ɽb5ǽ�cŽ��ý6�½P   P   9zýSýfvý��ý
�Ľ��Ž��ƽ��ǽcɽ�ɽx�ʽ��ʽ�ʽ�ʽeɽ�ǽb�ƽ��Ž�Ľ��ýP   P   KŽ?ŽS=Ž�EŽk[Ž�Ž�Žt$ƽ��ƽ��ƽ�Oǽ��ǽ^�ǽUǽǽ"�ƽT0ƽM�Ž��Ž�cŽP   P   ��ǽ��ǽ=Ƚ��ǽ��ǽ�*ǽ7�ƽ�#ƽ��Ž�iŽ�6Ž�Ž�Ž� Ž&>Ž�sŽ��ŽU0ƽb�ƽc5ǽP   P   �dʽ$I˽m�˽&�˽!C˽J[ʽ[*ɽ)�ǽݍƽ:hŽ5�Ľ�ýp�ýW�ýg�ý`�Ľ�sŽ"�ƽ�ǽ76ɽP   P   �>ͽ��ν�н�gнXнM�νz3ͽ(˽� ɽ��ƽ	4Ž'�ýý|�½"ýh�ý&>Žǽfɽ�4˽P   P   `�Ͻt�ҽ�wԽ�ս�սgqԽ�{ҽ��ϽF�̽N�ɽ�Iǽ�Ž��ý��½|�½W�ý� ŽUǽ�ʽ=�̽P   P   ҽ|�ս6�ؽ=�ڽ�?۽��ڽ��ؽ��սҽ�Bν!�ʽyxǽ�Ž��ýýp�ý�Ž_�ǽ �ʽ�OνP   P   h�ӽؽܽ�߽�����}߽
ܽxؽ%�ӽ��ν��ʽyxǽ�Ž'�ý�ý�Ž��ǽ��ʽ�ϽP   P   �Խ�XٽU޽�o��%�s潝!��h�?K޽yMٽ�Խ��ν!�ʽ�Iǽ	4Ž5�Ľ�6Ž�Oǽy�ʽ�ϽP   P   W�ӽ9Wٽ߽?佚轺*�U)�7�T7��߽yMٽ$�ӽ�BνM�ɽ��ƽ:hŽ�iŽ��ƽ�ɽ�JνP   P   ҽ�ؽ�R޽5>�3"�N]�~��Z�m�S7�?K޽xؽҽF�̽� ɽݍƽ��Ž��ƽcɽ��̽P   P   t�ϽH�սܽ�m�6轣]� ����Z�7��h�
ܽ��ս��Ͻ(˽)�ǽ�#ƽt$ƽ��ǽ+˽P   P   �4ͽF}ҽl�ؽ�߽}#�+�A~���~�T)꽜!�|߽��ؽ�{ҽy3ͽ[*ɽ7�ƽ�Ž��ƽ�*ɽP   P   �Zʽ{�ν�pԽ�ڽx����+꽢]�M]콺*�r���ཕ�ڽfqԽL�νJ[ʽ�*ǽ�Ž��Ž�*ǽP   P   [�ǽ1@˽��Ͻc|ս�;۽x��}#�5�2"齙��%��ཛ?۽�սWн!C˽��ǽj[Ž
�ĽOZŽP   P   �BŽ��ǽM�˽bнc|ս�ڽ�߽�m�4>�?��o⽔߽<�ڽ�ս�gн&�˽��ǽ�EŽ��ý@�ýP   P   �sý�8Ž�ȽM�˽��Ͻ�pԽl�ؽܽ�R޽߽U޽ܽ5�ؽ�wԽ�нl�˽<ȽS=Žfvý��½P   P   �R½>Oý�8Ž��ǽ1@˽{�νF}ҽG�ս�ؽ8Wٽ�Xٽؽ{�սs�ҽ��ν#I˽��ǽ?ŽSýFT½P   P   �RŽ}�Ž�xƽ��ǽs�ɽf�˽4�ͽ��Ͻeѽ�uҽ��ҽxҽjѽo�Ͻ/�ͽ_�˽k�ɽ��ǽ�}ƽ��ŽP   P   ��Žb�Ž�ƽ*�ƽ�ǽ�Jɽ��ʽ�I̽�ͽ��ν�Ͻ+ Ͻ��νP�ͽAQ̽��ʽ9Sɽ��ǽs�ƽRƽP   P   �}ƽ�_ƽ�zƽ��ƽFXǽ&Ƚ��Ƚ>�ɽ��ʽf˽D�˽�̽2�˽�k˽��ʽ�ɽ��ȽȽ�_ǽs�ƽP   P   ��ǽ��ǽ��ǽV�ǽ��ǽIȽ_EȽ)�Ƚ��Ƚ�#ɽ aɽŃɽ$�ɽ�eɽX*ɽ��Ƚ��Ƚ�NȽȽ��ǽP   P   l�ɽ5�ɽ��ɽ��ɽR�ɽ�Jɽ��Ƚs�Ƚp6Ƚ��ǽ�ǽS�ǽ��ǽ]�ǽ*�ǽe�ǽ�@Ƚ��Ƚ��Ƚ9SɽP   P   `�˽�\̽�̽)�̽$X̽��˽}�ʽ��ɽ��Ƚ��ǽUDǽ1�ƽ��ƽf�ƽ}�ƽ�Kǽe�ǽ��Ƚ�ɽ��ʽP   P   0�ͽuϽ��Ͻd$нi�Ͻ�Ͻ8�ͽTG̽��ʽ� ɽ��ǽ��ƽ�$ƽ1�Ž?(ƽ}�ƽ+�ǽX*ɽ��ʽBQ̽P   P   p�ϽQ�ѽY!ӽ`�ӽ��ӽ9ӽ��ѽu�Ͻ�ͽ~a˽�\ɽw�ǽ��ƽ��Ž1�Žf�ƽ]�ǽ�eɽ�k˽Q�ͽP   P   jѽrԽG,ֽ��׽�ؽM�׽�%ֽ�ӽ�_ѽ��νt�˽\}ɽ�ǽ��ƽ�$ƽ��ƽ��ǽ%�ɽ2�˽��νP   P    xҽI�ս��ؽP�ڽ5�۽l�۽��ڽ(�ؽ��ս�nҽ�Ͻ�̽\}ɽw�ǽ��ƽ1�ƽS�ǽŃɽ�̽, ϽP   P   ��ҽ$�ֽHڽ�7ݽ�%߽��߽~"߽Q2ݽS@ڽ��ֽ�ҽ�Ͻt�˽�\ɽ��ǽUDǽ�ǽ aɽD�˽�ϽP   P   �uҽ	�ֽ��ڽ��޽�=ὑ�����9��{޽<�ڽ��ֽ�nҽ��ν~a˽� ɽ��ǽ��ǽ�#ɽf˽��νP   P   eѽ�ս!Fڽ��޽t���>��	��<�����{޽S@ڽ��ս�_ѽ�ͽ��ʽ��Ƚp6Ƚ��Ƚ��ʽ�ͽP   P   ��Ͻ�Խģؽ�5ݽ�<�
?�P��`���<��9�Q2ݽ(�ؽ�ӽt�ϽTG̽��ɽr�Ƚ*�Ƚ>�ɽ�I̽P   P   4�ͽخѽL'ֽA�ڽ�#߽���
�P���	���~"߽��ڽ�%ֽ��ѽ7�ͽ}�ʽ�Ƚ_EȽ��Ƚ �ʽP   P   f�˽iϽ�ӽ��׽�۽��߽���
?��>佐����߽l�۽L�׽8ӽ�Ͻ��˽�JɽIȽ&Ƚ�JɽP   P   t�ɽ�U̽��Ͻ�ӽؽ�۽�#߽�<�t���=Ὥ%߽4�۽�ؽ��ӽi�Ͻ$X̽R�ɽ��ǽFXǽ�ǽP   P   ��ǽ �ɽy�̽�н�ӽ��׽A�ڽ�5ݽ��޽��޽�7ݽO�ڽ��׽`�ӽc$н)�̽��ɽV�ǽ��ƽ*�ƽP   P   �xƽ�ǽ]�ɽy�̽��Ͻ�ӽK'ֽãؽ!Fڽ��ڽHڽ��ؽF,ֽX!ӽ��Ͻ�̽��ɽ��ǽ�zƽ�ƽP   P   }�Ž�\ƽ�ǽ �ɽ�U̽iϽ׮ѽ�Խ�ս�ֽ#�ֽI�սqԽP�ѽuϽ�\̽5�ɽ��ǽ�_ƽb�ŽP   P   x�ǽAȽ�Ƚ��ɽ� ˽ �̽�:ν	�Ͻ��нO�ѽ��ѽ��ѽ��н�Ͻ�@ν��̽�&˽��ɽ��Ƚ-ȽP   P   -Ƚ�Ƚ�iȽ\ɽE�ɽ��ʽ�̽�ͽ�νN�ν�2Ͻ�3Ͻ}�ν�ν�#ͽ�	̽��ʽ��ɽrɽ�lȽP   P   ��Ƚ�Ƚb�ȽɽLlɽ��ɽ��ʽ6H˽B�˽s̽�̽,�̽��̽]w̽j�˽HO˽{�ʽ$�ɽrɽrɽP   P   ��ɽ��ɽ��ɽ�ɽ��ɽ�ɽ1!ʽTʽO�ʽ^�ʽ��ʽ�	˽�
˽��ʽ��ʽW�ʽ�[ʽ�(ʽ$�ɽ��ɽP   P   �&˽�O˽]˽�L˽?"˽�ʽ��ʽ�Sʽ*ʽ�ɽ��ɽF�ɽܪɽ��ɽ��ɽz�ɽʽ�[ʽ{�ʽ��ʽP   P   ��̽?)ͽ]jͽiͽP%ͽg�̽n̽G˽?�ʽ>�ɽrZɽ��Ƚ��ȽS�Ƚ5�Ƚ`ɽz�ɽW�ʽHO˽�	̽P   P   �@ν)Ͻ�Ͻ��ϽW�Ͻ$Ͻ�9ν�ͽ��˽��ʽ��ɽ��Ƚ�Ƚ�VȽC�Ƚ5�Ƚ��ɽ��ʽk�˽�#ͽP   P   �Ͻ�ѽ'ҽZ�ҽҲҽ #ҽ�ѽ��Ͻ�ν>o̽��ʽ�ɽ��Ƚ�UȽ�VȽS�Ƚ��ɽ��ʽ]w̽�νP   P   ��нa�ҽ�_Խ�bս�սj`ս}ZԽ��ҽ��н��ν��̽�˽a�ɽ��Ƚ�Ƚ��Ƚܪɽ�
˽��̽}�νP   P   ��ѽ{Խ-ֽú׽��ؽ�ؽ
�׽�'ֽ�Խ
�ѽ�,Ͻ��̽�˽�ɽ��Ƚ��ȽF�ɽ�	˽-�̽�3ϽP   P   ��ѽ��Խ�Y׽�wٽ�ڽ�S۽��ڽ�sٽ�S׽<�Խ��ѽ�,Ͻ��̽��ʽ��ɽrZɽ��ɽ��ʽ�̽�2ϽP   P   O�ѽɽԽ��׽�dڽXܽ�aݽ�`ݽ(UܽY`ڽ�׽<�Խ
�ѽ��ν>o̽��ʽ>�ɽ�ɽ^�ʽs̽O�νP   P   ��н�ԽX׽�cڽB�ܽLz޽�	߽�x޽��ܽY`ڽ�S׽�Խ��н�ν��˽?�ʽ*ʽO�ʽB�˽�νP   P   	�ϽI�ҽ+*ֽrvٽ�WܽSz޽1�߽߽͝�x޽(Uܽ�sٽ�'ֽ��ҽ��Ͻ�ͽG˽�SʽTʽ6H˽�ͽP   P   �:ν�ѽ\Խ\�׽��ڽ�aݽ>
߽1�߽�	߽�`ݽ��ڽ	�׽|ZԽ�ѽ�9νm̽��ʽ1!ʽ��ʽ�̽P   P    �̽�#Ͻ�"ҽ�_սӌؽ�S۽�aݽRz޽Kz޽�aݽ�S۽�ؽj`ս�"ҽ$Ͻg�̽�ʽ�ɽ��ɽ��ʽP   P   � ˽�#ͽ��Ͻ��ҽO�սӌؽ��ڽ�WܽA�ܽXܽ�ڽ��ؽ�սҲҽW�ϽP%ͽ>"˽��ɽLlɽE�ɽP   P   ��ɽ�J˽+fͽ��Ͻ��ҽ�_ս[�׽rvٽ�cڽ�dڽ�wٽú׽�bսZ�ҽ��Ͻiͽ�L˽�ɽɽ\ɽP   P   �Ƚ��ɽ5Y˽+fͽ��Ͻ�"ҽ\Խ**ֽX׽��׽Y׽-ֽ�_Խ'ҽ�Ͻ]jͽ]˽��ɽb�Ƚ�iȽP   P   AȽo�Ƚ��ɽ�J˽�#ͽ�#Ͻ�ѽH�ҽ�ԽȽԽ��Խ{Խa�ҽ�ѽ)Ͻ?)ͽ�O˽��ɽ�Ƚ�ȽP   P   ��ɽ��ɽxʽ�?˽�@̽]dͽ�ν��ϽY�нlѽ(GѽDѽ�нU�Ͻ��ν�iͽ�D̽�C˽C{ʽ��ɽP   P   ��ɽ��ɽ�7ʽ�ʽ�N˽�̽�̽�ͽ#sν��ν�DϽEϽX�νLwν(�ͽ^�̽̽T˽��ʽu:ʽP   P   C{ʽ�hʽ�yʽg�ʽ}�ʽde˽H�˽�`̽�̽H<ͽ�}ͽ��ͽ�ͽ�?ͽ��̽qf̽�˽*k˽� ˽��ʽP   P   �C˽�;˽�:˽A˽AO˽ye˽��˽�˽�˽��˽�̽,̽;-̽r̽P ̽��˽g�˽�˽*k˽T˽P   P   �D̽=b̽)l̽&`̽@A̽�̽��˽ɪ˽V{˽�T˽�:˽�*˽�%˽�,˽J>˽Z˽�˽g�˽�˽̽P   P   �iͽw�ͽ��ͽA�ͽ�ͽ�dͽo�̽�_̽�˽T˽��ʽ%�ʽ�~ʽ	�ʽm�ʽ��ʽZ˽��˽qf̽^�̽P   P   ��ν>Ͻ=�Ͻ7�Ͻ8�ϽF:ϽA�ν��ͽ?�̽
�˽9˽��ʽQEʽ%ʽ�Fʽm�ʽJ>˽P ̽��̽(�ͽP   P   U�Ͻ�н}pѽ��ѽt�ѽ[mѽ4�н��Ͻ�pν*9ͽ�̽'(˽ }ʽ�#ʽ%ʽ	�ʽ�,˽r̽�?ͽLwνP   P   �н��ѽ2ӽ��ӽ2Խ��ӽuӽ`�ѽ0н�νzͽ(̽�"˽ }ʽQEʽ�~ʽ�%˽<-̽�ͽY�νP   P   Dѽ��ҽH`Խ́սPֽֽ�~ս`\Խe�ҽ�ѽ�?Ͻ��ͽ(̽'(˽��ʽ%�ʽ�*˽,̽��ͽEϽP   P   (GѽPUӽ�:սL�ֽ;�׽�ؽ�׽�ֽe6ս^Pӽ�Aѽ�?Ͻzͽ�̽9˽��ʽ�:˽�̽�}ͽ�DϽP   P   lѽ�Tӽ�ս_m׽��ؽ�ٽ"�ٽ{�ؽ3j׽�ս^Pӽ�ѽ�ν*9ͽ
�˽T˽�T˽��˽I<ͽ��νP   P   Y�н��ҽ�9ս
m׽�4ٽ�]ڽ�ڽP\ڽ�2ٽ3j׽e6սe�ҽ0н�pν?�̽�˽V{˽�˽�̽#sνP   P   ��Ͻ>�ѽG^Խ��ֽU�ؽ>]ڽt-۽n-۽P\ڽ{�ؽ�ֽ_\Խ`�ѽ��Ͻ��ͽ�_̽ɪ˽�˽�`̽�ͽP   P   �ν�н�ӽ�ս��׽��ٽ��ڽt-۽�ڽ"�ٽ�׽�~սuӽ3�н@�νo�̽��˽��˽H�˽�̽P   P   ]dͽ�9Ͻ�lѽH�ӽ�ֽ�ؽ��ٽ>]ڽ�]ڽ�ٽ�ؽֽ��ӽZmѽF:Ͻ�dͽ�̽ye˽de˽�̽P   P   �@̽�ͽԨϽ'�ѽԽ�ֽ��׽U�ؽ�4ٽ��ؽ;�׽Oֽ2Խt�ѽ8�Ͻ�ͽ@A̽AO˽}�ʽ�N˽P   P   �?˽A^̽��ͽ��Ͻ'�ѽH�ӽ�ս��ֽ
m׽^m׽L�ֽˁս��ӽ��ѽ7�ϽA�ͽ&`̽A˽g�ʽ�ʽP   P   xʽ�8˽�i̽��ͽԨϽ�lѽ�ӽG^Խ�9ս�ս�:սG`Խ1ӽ}pѽ=�Ͻ��ͽ(l̽�:˽�yʽ�7ʽP   P   ��ɽgʽ�8˽A^̽�ͽ�9Ͻ �н>�ѽ��ҽ�TӽOUӽ��ҽ��ѽ�н>Ͻw�ͽ=b̽�;˽�hʽ��ɽP   P   �A˽Ib˽w�˽)W̽mͽ�ͽ�νG�Ͻ�<нϧн��н8�н�>н�Ͻ��ν7�ͽ�ͽPZ̽��˽rc˽P   P   rc˽�b˽��˽��˽�b̽~�̽̕ͽ�1νM�ν=ϽLRϽ�RϽWϽ��ν�5ν�ͽ��̽�f̽��˽�˽P   P   ��˽z�˽E�˽��˽<%̽iu̽��̽//ͽ��ͽ��ͽnν�ν�ν}�ͽ�ͽ�3ͽc�̽�y̽�(̽��˽P   P   PZ̽T̽�R̽%X̽�b̽�u̽B�̽_�̽��̽�̽x�̽ͽͽ��̽��̽U�̽��̽�̽�y̽�f̽P   P   �ͽy/ͽ}5ͽ�-ͽ�ͽ��̽��̽_�̽�̽�g̽�R̽�E̽�B̽XG̽�U̽l̽m�̽��̽c�̽��̽P   P   7�ͽ�5ν�Wν(Wν�2ν�ͽR�ͽ�.ͽ��̽!g̽{̽��˽t�˽;�˽��˽�̽l̽U�̽�3ͽ�ͽP   P   ��ν|MϽ��ϽɺϽ�Ͻ�JϽl�ν�0νF�ͽ��̽�Q̽��˽�˽��˽�˽��˽�U̽��̽�ͽ�5νP   P   �Ͻ]н!�н#7ѽ6ѽ��нYнޗϽ`�ν]�ͽ>�̽�C̽��˽f�˽��˽;�˽XG̽��̽}�ͽ��νP   P   �>н�GѽEҽĦҽ��ҽ]�ҽ�ҽ`Cѽ2:нdϽ��ͽ	ͽl@̽��˽�˽t�˽�B̽ͽ�νWϽP   P   8�н�ѽZӽM�ӽ/SԽmRԽ��ӽRӽ��ѽפнbNϽ�ν	ͽ�C̽��˽��˽�E̽ͽ�ν�RϽP   P   ��нGOҽ!�ӽ��Խ�ս?�ս��ս��Խ
�ӽbKҽ��нaNϽ��ͽ>�̽�Q̽{̽�R̽x�̽nνLRϽP   P   ϧн�Nҽ��ӽ�HսKMֽ��ֽ��ֽ�KֽsFս��ӽbKҽפнdϽ]�ͽ��̽!g̽�g̽�̽��ͽ=ϽP   P   �<н��ѽ5�ӽ�Hսˑֽ�g׽�׽�f׽;�ֽsFս
�ӽ��ѽ1:н`�νF�ͽ��̽�̽��̽��ͽM�νP   P   G�Ͻ�Dѽ�ӽa�Խ-Mֽ�g׽��׽��׽�f׽�Kֽ��ԽRӽ`CѽޗϽ�0ν�.ͽ_�̽_�̽//ͽ�1νP   P   �ν�YнYҽ��ӽl�սS�ֽı׽��׽�׽��ֽ��ս��ӽ�ҽYнl�νQ�ͽ��̽B�̽��̽̕ͽP   P   �ͽ?JϽ��н��ҽ3RԽK�սS�ֽ�g׽�g׽��ֽ?�սmRԽ]�ҽ��н�JϽ~�ͽ��̽�u̽iu̽~�̽P   P   mͽM2ν�Ͻ5ѽ��ҽ3RԽl�ս-MֽʑֽKMֽ�ս/SԽ��ҽ6ѽ�Ͻ�2ν�ͽ�b̽<%̽�b̽P   P   )W̽9,ͽ6UνظϽ5ѽ��ҽ��ӽa�Խ�Hս�Hս��ԽM�ӽĦҽ"7ѽɺϽ(Wν�-ͽ%X̽��˽��˽P   P   w�˽`Q̽�3ͽ6Uν�Ͻ��нYҽ�ӽ5�ӽ��ӽ!�ӽZӽEҽ �н��Ͻ�Wν}5ͽ�R̽E�˽��˽P   P   Ib˽�˽`Q̽9,ͽM2ν?JϽ�Yн�Dѽ��ѽ�NҽGOҽ�ѽ�Gѽ]н|MϽ�5νx/ͽT̽y�˽�b˽P   P   Y̽�o̽��̽�&ͽG�ͽ�Wν1�ν�Ͻ�	нYн�sн�Yн�нe�Ͻ�ν�Zν �ͽ+)ͽ+�̽�p̽P   P   �p̽�o̽�̽��̽�/ͽd�ͽ�ν@�ν��νB5Ͻt\ϽC]Ͻ�6Ͻz�νq�ν�ν�ͽ�2ͽ��̽��̽P   P   +�̽{�̽W�̽��̽&ͽ�=ͽ�ͽ��ͽ�ν�@ν1cνapν)dν�Bνfν>�ͽ��ͽyAͽͽ��̽P   P   +)ͽ�#ͽ�"ͽ?'ͽ40ͽ�=ͽuOͽ?eͽ�{ͽ�ͽ:�ͽ?�ͽשͽ@�ͽ��ͽ@ͽ1iͽGSͽyAͽ�2ͽP   P   �ͽ��ͽ��ͽ��ͽ��ͽ��ͽςͽ+eͽPJͽ�3ͽM#ͽ�ͽaͽ�ͽV%ͽ!7ͽ�Mͽ1iͽ��ͽ�ͽP   P   �ZνF�ν��ν6�ν4�ν�Wν*ν/�ͽ{ͽq3ͽ\�̽�̽��̽Y�̽�̽e�̽!7ͽ@ͽ?�ͽ�νP   P   �νCZϽ��Ͻ�ϽY�ϽXϽ��ν�νj
ν �ͽI"ͽ��̽0�̽�̽M�̽�̽V%ͽ��ͽfνq�νP   P   e�Ͻ�"н��н��н�н��н�н��Ͻw�ν�>ν��ͽ�ͽ��̽G�̽�̽Y�̽�ͽ@�ͽ�Bν{�νP   P   �н
�нkѽ��ѽ��ѽ?�ѽ�hѽ�н�н3Ͻ�`ν�ͽ3ͽ��̽0�̽��̽aͽשͽ)dν�6ϽP   P   �Yн�Lѽ�ҽ��ҽ�ӽ`ӽ�ҽ2ҽ�Iѽ�Vн�YϽ6mν�ͽ�ͽ��̽�̽�ͽ?�ͽbpνD]ϽP   P   �sн͎ѽؑҽFbӽT�ӽ=ԽH�ӽF`ӽ��ҽ�ѽ�pн�YϽ�`ν��ͽI"ͽ\�̽M#ͽ:�ͽ1cνt\ϽP   P   Yн��ѽ��ҽR�ӽlyԽa�Խ��Խ�xԽm�ӽ
�ҽ�ѽ�Vн3Ͻ�>ν �ͽq3ͽ�3ͽ�ͽ�@νB5ϽP   P   �	н�Kѽ:�ҽ�ӽ{�Խ;Eս�zս�Dս(�Խm�ӽ��ҽ�Iѽ�нv�νj
ν{ͽPJͽ�{ͽ�ν��νP   P   �Ͻ�н�ҽ�aӽ>yԽ=Eս��ս��ս�Dս�xԽF`ӽ2ҽ�н��Ͻ�ν/�ͽ+eͽ?eͽ��ͽ@�νP   P   1�νS нsiѽT�ҽ��ӽ)�ԽF{ս��ս�zս��ԽH�ӽ�ҽ�hѽ�н��ν*νςͽuOͽ�ͽ�νP   P   �Wν�WϽ��нG�ѽ%ӽ=Խ)�Խ=Eս;Eսa�Խ=Խ`ӽ?�ѽ��нXϽ�Wν��ͽ�=ͽ�=ͽd�ͽP   P   G�ͽ��ν��Ͻ�н1�ѽ%ӽ��ӽ=yԽ{�ԽlyԽT�ӽ�ӽ��ѽ�нY�Ͻ4�ν��ͽ40ͽ&ͽ�/ͽP   P   �&ͽ]�ͽޡν��Ͻ�нG�ѽT�ҽ�aӽ�ӽR�ӽFbӽ��ҽ��ѽ��н�Ͻ6�ν��ͽ?'ͽ��̽��̽P   P   ��̽�!ͽ�ͽޡν��Ͻ��нsiѽ�ҽ:�ҽ��ҽؑҽ�ҽkѽ��н��Ͻ��ν��ͽ�"ͽW�̽�̽P   P   �o̽�̽�!ͽ]�ͽ��ν�WϽS н�н�Kѽ��ѽ͎ѽ�Lѽ
�н�"нCZϽF�ν��ͽ�#ͽ{�̽�o̽P   P   �%ͽA8ͽ�mͽ)�ͽO+ν��ν�Ͻ��Ͻ3�Ͻ�н;3н0н��Ͻ��ϽRϽإν�-ν2�ͽoͽ�8ͽP   P   �8ͽC8ͽGRͽ�ͽ��ͽ.νdrν��ν�Ͻ_HϽ�dϽpeϽ|IϽ�Ͻ�νuν�ν��ͽ.�ͽ�SͽP   P   oͽ5gͽanͽ��ͽ�ͽ��ͽ"ν ;ν�jν��νܬνP�ν��ν=�ν\mν�=ν:	ν��ͽ��ͽ.�ͽP   P   2�ͽ��ͽr�ͽi�ͽ��ͽ��ͽ��ͽ��ͽν�νLν}!ν�!ν�ν�ν�νl�ͽ��ͽ��ͽ��ͽP   P   �-ν�8ν`<ν�7ν�+νIν#νU�ͽ(�ͽ��ͽ��ͽ��ͽ��ͽ��ͽS�ͽ3�ͽ{�ͽl�ͽ:	ν�νP   P   إνd�ν��ν��ν�νq�ν'rν�:ν� ν��ͽA�ͽ�ͽ�nͽooͽ��ͽ֠ͽ3�ͽ�ν�=νuνP   P   RϽ�cϽ��Ͻ��Ͻ�Ͻ�aϽ�Ͻ4�ν�iν�ν��ͽ�~ͽ�Vͽ�Hͽ�Wͽ��ͽS�ͽ�ν\mν�νP   P   ��Ͻ~�Ͻ�Cн7lнlн)BнG�Ͻ��Ͻ�Ͻ[�ν�ν��ͽnͽ�Hͽ�Hͽooͽ��ͽ�ν=�ν�ϽP   P   ��Ͻ%uнG�н�2ѽLѽ�1ѽ��н�rн��Ͻ�FϽ��ν�νu�ͽnͽ�Vͽ�nͽ��ͽ�!ν��ν|IϽP   P   0нJ�н�kѽV�ѽ|ҽ2ҽ]�ѽ�iѽ��н�н�bϽӳν�ν��ͽ�~ͽ�ͽ��ͽ}!νP�νpeϽP   P   ;3н!ѽT�ѽ�XҽȺҽ��ҽǹҽ7Wҽ��ѽ�ѽ�0н�bϽ��ν�ν��ͽA�ͽ��ͽLνܬν�dϽP   P   �н�ѽ��ѽl�ҽ�#ӽmӽ�lӽ�"ӽ��ҽ��ѽ�ѽ�н�FϽ[�ν�ν��ͽ��ͽ�ν��ν`HϽP   P   3�Ͻ��н��ѽ�ҽsHӽa�ӽ��ӽ�ӽWGӽ��ҽ��ѽ��н��Ͻ�Ͻ�iν� ν(�ͽν�jν�ϽP   P   ��Ͻtн�jѽXҽO#ӽ��ӽYԽ&Խ�ӽ�"ӽ7Wҽ�iѽ�rн��Ͻ4�ν�:νU�ͽ��ͽ ;ν��νP   P   �Ͻ��Ͻ��н`�ѽ��ҽmӽ��ӽYԽ��ӽ�lӽǹҽ]�ѽ��нG�Ͻ�Ͻ'rν#ν��ͽ"νdrνP   P   ��ν�aϽ)Bн�1ѽ	ҽ��ҽmӽ��ӽa�ӽmӽ��ҽ2ҽ�1ѽ)Bн�aϽq�νIν��ͽ��ͽ.νP   P   O+ν��νJ�Ͻ*kнeKѽ	ҽ��ҽO#ӽsHӽ�#ӽǺҽ|ҽLѽlн�Ͻ�ν�+ν��ͽ�ͽ��ͽP   P   )�ͽ7ν��ν��Ͻ*kн�1ѽ`�ѽXҽ�ҽl�ҽ�XҽV�ѽ�2ѽ7lн��Ͻ��ν�7νi�ͽ��ͽ�ͽP   P   �mͽ��ͽ;ν��νJ�Ͻ)Bн��н�jѽ��ѽ��ѽS�ѽ�kѽG�н�Cн��Ͻ��ν`<νr�ͽanͽGRͽP   P   A8ͽ fͽ��ͽ7ν��ν�aϽ��Ͻtн��н�ѽ!ѽJ�н%uн~�Ͻ�cϽd�ν�8ν��ͽ4gͽC8ͽP   P   ��ͽJ�ͽ��ͽK4ν��ν5�ν#6Ͻs�Ͻ��Ͻ��Ͻ�н��Ͻ�Ͻ!�Ͻ8Ͻ��ν�ν�5ν��ͽ��ͽP   P   ��ͽ��ͽu�ͽ�νA:ν�wν�ν�νw-ϽUϽ0jϽ�jϽ
VϽ�.Ͻ��ν�ν�yν�;νEνe�ͽP   P   ��ͽ��ͽ��ͽν ν�Aνygν��νf�ν[�ν��νS�νA�ν��ν��νːν�iν�CνG"νEνP   P   �5νD2ν�1ν�4νE:ν�Aν�Kν�Wν�cνgoν�vν�{ν�{νxν�pν�eν�YνKNν�Cν�;νP   P   �ν��νv�ν�ν&�ν�wν�gνJWν�Gν�;ν�1ν�+ν+ν�,νH3ν�=ν�Jν�Yν�iν�yνP   P   ��ν��ν�Ͻ�Ͻ!�ν2�ν��ν[�ν�cν�;ννUν�ͽF�ͽνν�=ν�eνːν�νP   P   8Ͻ�iϽA�Ͻ��ϽK�Ͻ�gϽ6Ͻk�νʱνjnν.1ν�ν��ͽ��ͽ��ͽνH3ν�pν��ν��νP   P   "�Ͻ��Ͻ^н�,н�,н=н6�Ͻ͇Ͻ_,Ͻ��ν�uνc+νO�ͽ��ͽ��ͽF�ͽ�,νxν��ν�.ϽP   P   �Ͻ�4н��нP�н��нF�нb�н�2н��Ͻ�SϽ��νOzν�)νO�ͽ��ͽ�ͽ+ν�{νA�ν
VϽP   P   ��Ͻ�xнa�н�;ѽ|fѽ9fѽG;ѽ��н�vн��Ͻ�hϽm�νOzνc+ν�νUν�+ν�{νS�ν�jϽP   P   �н�н�'ѽz�ѽR�ѽ��ѽ��ѽi�ѽ�&ѽ�нн�hϽ��ν�uν.1νν�1ν�vν��ν0jϽP   P   ��Ͻu�н�<ѽm�ѽ4,ҽ�`ҽ�`ҽ{+ҽd�ѽ;ѽ�н��Ͻ�SϽ��νjnν�;ν�;νgoν[�νUϽP   P   ��Ͻ�wн�'ѽi�ѽ�Fҽ#�ҽ�ҽ�ҽGFҽd�ѽ�&ѽ�vн��Ͻ_,Ͻʱν�cν�Gν�cνf�νw-ϽP   P   s�Ͻ�3н��н��ѽ�+ҽ4�ҽ!�ҽ��ҽ�ҽ{+ҽi�ѽ��н�2н̇Ͻk�ν[�νJWν�Wν��ν�νP   P   #6Ͻ��Ͻb�нZ;ѽ3�ѽaҽ��ҽ!�ҽ�ҽ�`ҽ��ѽG;ѽa�н6�Ͻ6Ͻ��ν�gν�Kνygν�νP   P   5�ν&hϽ=н��н=fѽ�ѽaҽ4�ҽ#�ҽ�`ҽ��ѽ9fѽF�н=н�gϽ2�ν�wν�Aν�Aν�wνP   P   ��ν��ν��Ͻ�+н��н=fѽ3�ѽ�+ҽ�Fҽ4,ҽR�ѽ|fѽ��н�,нK�Ͻ!�ν&�νE:ν νA:νP   P   K4ν��νPϽ�Ͻ�+н��нZ;ѽ��ѽi�ѽm�ѽy�ѽ�;ѽP�н�,н��Ͻ�Ͻ�ν�4νν�νP   P   ��ͽ71νH�νPϽ��Ͻ=нa�н��н�'ѽ�<ѽ�'ѽa�н��н^н@�Ͻ�Ͻv�ν�1ν��ͽu�ͽP   P   J�ͽ��ͽ71ν��ν��ν&hϽ��Ͻ�3н�wнu�н�н�xн�4н��Ͻ�iϽ��ν��νD2ν��ͽ��ͽP   P   �3νx=ν�Zν�ν��ν�Ͻ�GϽ(�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻl�ϽdIϽ$Ͻ8�ν �ν�[ν�=νP   P   �=ν>νGLν{hνs�νz�ν��ν	ϽsBϽ0`Ͻ�oϽpϽ�`Ͻ?CϽaϽ�ν��ν��νxiν"MνP   P   �[ν�Vν�Zν�hν@{ν��ν��ν��νq�ν��ν�
ϽXϽ9Ͻ��ν&�ν��νY�ν��ν�|νxiνP   P    �νD�ν	�ν��νT�ν,�ν@�ν�νc�ν�ν$�νV�ν��νĻν+�νԮνʦν
�ν��ν��νP   P   8�νZ�ν��ν��ν��νv�νy�ν��ν��ν׎ν�νN�νt�ν�νM�ν�ν��νʦνY�ν��νP   P   $Ͻ�Ͻ%Ͻ�$Ͻ�Ͻ�Ͻ.�ν��ν�νێν
wνteν�[ν�[νAfνVxν�νԮν��ν�νP   P   eIϽoϽ̆Ͻ��Ͻ2�Ͻ�mϽ�GϽ�Ͻ�ν4�ν͇νeν+NνEFν�NνAfνM�ν,�ν&�νaϽP   P   l�Ͻp�Ͻ��Ͻ��Ͻ��Ͻ��ϽB�Ͻ��ϽcAϽ4�ν-�ν��ν3[νFνEFν�[ν�νĻν��ν@CϽP   P   ��Ͻ�н*Bн	jнxxнOiн3AнVнl�Ͻ_Ͻ�	Ͻ3�νd�ν3[ν+Nν�[νt�ν��ν9Ͻ�`ϽP   P   ��ϽU6нd�н��нU�н�н��н-�н5н5�ϽlnϽϽ3�ν��νeνteνN�νV�νXϽpϽP   P   ��ϽQнG�н�ѽ�=ѽ�Oѽ
=ѽ�ѽ6�нwOнt�ϽlnϽ�	Ͻ-�ν͇ν
wν�ν$�ν�
Ͻ�oϽP   P   ��Ͻ�Pн��н,ѽ!vѽ��ѽ}�ѽvuѽg+ѽ��нwOн5�Ͻ_Ͻ4�ν4�νێν׎ν�ν��ν0`ϽP   P   �Ͻ�5н��нC,ѽK�ѽX�ѽW�ѽ�ѽÈѽg+ѽ6�н5нl�ϽbAϽ�ν�ν��νc�νr�νsBϽP   P   (�Ͻ8н�нѽ�uѽ�ѽ��ѽJ�ѽ�ѽvuѽ�ѽ-�нVн��Ͻ�Ͻ��ν��ν�ν��ν	ϽP   P   �GϽ��ϽAн<�нC=ѽȜѽT�ѽ��ѽW�ѽ}�ѽ
=ѽ��н3AнB�Ͻ�GϽ.�νy�ν@�ν��ν��νP   P   �Ͻ�mϽ��Ͻ�iн?�нbOѽȜѽ�ѽX�ѽ��ѽ�Oѽ�нOiн��Ͻ�mϽ�Ͻv�ν,�ν��νz�νP   P   ��ν�Ͻ{�ϽI�Ͻ�wн?�нC=ѽ�uѽK�ѽ!vѽ�=ѽT�нxxн��Ͻ2�Ͻ�Ͻ��νT�ν@{νs�νP   P   �νt�ν$Ͻq�ϽI�Ͻ�iн<�нѽC,ѽ,ѽ�ѽ��н	jн��Ͻ��Ͻ�$Ͻ��ν��ν�hν{hνP   P   �Zνn�ν��ν$Ͻ{�Ͻ��ϽAн�н��н��нG�нd�н*Bн��Ͻ̆Ͻ%Ͻ��ν�ν�ZνGLνP   P   x=ν�Vνn�νt�ν�Ͻ�mϽ��Ͻ8н�5н�PнQнU6н�нp�ϽoϽ�ϽZ�νD�ν�Vν>νP   P   ��ν�ν��ν��νT�ν�%ϽWϽكϽ�Ͻk�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ2XϽ'ϽK�νU�νԧνA�νP   P   A�νm�νܚν¯νm�ν��νϽ�4Ͻ�RϽwgϽ�rϽ�rϽhϽfSϽ�5ϽϽM�ν��ν{�νj�νP   P   ԧν��ν�ν��νz�νl�ν��ν>�ν�ϽϽ�(Ͻ�,Ͻ&)Ͻ�Ͻ�Ͻ��νP�ν��ν��ν{�νP   P   U�ν��ν��ν�νv�ν��ν��ν��ν��νC�νM�νp�ν��ν��ν[�ν��ν-�ν��ν��ν��νP   P   K�ν��ν��ν7�νT�ν&�ν��ν��ν�ν��ν|�ν��νg�ν�νP�ν��νV�ν-�νP�νM�νP   P   'Ͻ�4Ͻ�;Ͻe;Ͻ=4Ͻ)&Ͻ�Ͻ;�νj�ν��ν��νݬν%�νF�ν��νi�ν��ν��ν��νϽP   P   2XϽ&sϽ�ϽʉϽt�ϽrϽ�VϽ�4Ͻ_Ͻ��ν�ν��ν�νa�νc�ν��νP�ν[�ν�Ͻ�5ϽP   P   ��Ͻk�Ͻ��Ͻ��Ͻ��Ͻ0�Ͻ��Ͻu�Ͻ�QϽ�Ͻ��ν�ν��ν�νa�νF�ν�ν��ν�ϽfSϽP   P   ��Ͻ�Ͻ�н�+н�5нe+нн��Ͻ��Ͻ�fϽ�'Ͻ��ν��ν��ν�ν%�νg�ν��ν&)ϽhϽP   P   �Ͻ�нvCн�oн��н�нMoн�Bн�н��Ͻ�qϽ�+Ͻ��ν�ν��νݬν��νp�ν�,Ͻ�rϽP   P   ��ϽLн�dн��н=�н:�н��н?�н�cн0н��Ͻ�qϽ�'Ͻ��ν�ν��ν|�νM�ν�(Ͻ�rϽP   P   k�Ͻ,н"qн��нc�нѽѽ	�н��нSpн0н��Ͻ�fϽ�Ͻ��ν��ν��νC�νϽwgϽP   P   �ϽYнldн��нv�н�+ѽ�:ѽ�+ѽ�н��н�cн�н��Ͻ�QϽ_Ͻj�ν�ν��ν�Ͻ�RϽP   P   كϽ6�ϽCн��нv�н�+ѽmIѽIIѽ�+ѽ	�н?�н�Bн��Ͻu�Ͻ�4Ͻ;�ν��ν��ν>�ν�4ϽP   P   WϽ��Ͻ/н�oн��н<ѽ�:ѽmIѽ�:ѽѽ��нMoнн��Ͻ�VϽ�Ͻ��ν��ν��νϽP   P   �%Ͻ7rϽ!�ϽD+нz�н@�н<ѽ�+ѽ�+ѽѽ:�н�нe+н0�ϽrϽ)&Ͻ&�ν��νl�ν��νP   P   T�ν�3Ͻ%�Ͻ~�Ͻn5нz�н��нv�нv�нc�н=�н��н�5н��Ͻt�Ͻ=4ϽT�νv�νz�νm�νP   P   ��ν��ν�:Ͻ=�Ͻ~�ϽD+н�oн��н��н��н��н�oн�+н��ϽʉϽe;Ͻ7�ν�ν��ν¯νP   P   ��ν7�νL�ν�:Ͻ%�Ͻ!�Ͻ/нCнldн"qн�dнvCн�н��Ͻ�Ͻ�;Ͻ��ν��ν�νܚνP   P   �ν~�ν7�ν��ν�3Ͻ7rϽ��Ͻ6�ϽYн,нLн�н�Ͻk�Ͻ&sϽ�4Ͻ��ν��ν��νm�νP   P   �ν�νR�ν��ν3Ͻ�<Ͻ;aϽ:�ϽۜϽ��ϽY�Ͻ��Ͻ�ϽłϽ�aϽ�=Ͻ�Ͻ|�ν��νk�νP   P   k�ν:�νs�ν�νg�ν�Ͻ�.ϽiGϽ9]Ͻ�mϽ<wϽHwϽ�mϽ2^Ͻ�HϽ�/Ͻ�Ͻv�ν��ν��νP   P   ��ν��νu�ν6�ν�ν��ν�ϽeϽq,Ͻ18Ͻm?Ͻ"BϽ�?Ͻ�8Ͻ�,ϽbϽ�Ͻ��ν��ν��νP   P   |�ν��ν��ν	�ν��ν��νϽϽ�Ͻ�Ͻ�ϽdϽ�Ͻ)Ͻ�Ͻ�Ͻ>	ϽAϽ��νv�νP   P   �Ͻ�ϽϽ=ϽϽϽ�ϽCϽVϽL�ν9�ν��ν �ν��ν��ν>�ν0Ͻ>	Ͻ�Ͻ�ϽP   P   �=Ͻ=HϽ3NϽ'NϽ�GϽ�<Ͻ�.Ͻ0ϽnϽ8�ν��ν��νO�ν��νR�ν>�ν>�ν�ϽbϽ�/ϽP   P   �aϽluϽ@�Ͻ��Ͻ�Ͻ�tϽ�`Ͻ_GϽ�+Ͻ�Ͻ��ν��ν��ν��ν��νR�ν��ν�Ͻ�,Ͻ�HϽP   P   łϽp�Ͻ��Ͻ��ϽL�Ͻ��ϽŠϽׁϽ�\Ͻ�7Ͻ=Ͻ@�ν�ν[�ν��ν��ν��ν)Ͻ�8Ͻ2^ϽP   P   �Ͻi�Ͻ��Ͻ��Ͻxн��Ͻ��Ͻt�Ͻ�Ͻ>mϽ�>Ͻ�ϽJ�ν�ν��νO�ν �ν�Ͻ�?Ͻ�mϽP   P   ��Ͻ��ϽIн|0н�Aн�Aн�/н�н�Ͻh�Ͻ\vϽGAϽ�Ͻ@�ν��ν��ν��νdϽ"BϽHwϽP   P   Y�Ͻ��Ͻ(н�Tн�pн�zн�pнPTн'нE�Ͻz�Ͻ\vϽ�>Ͻ=Ͻ��ν��ν9�ν�Ͻm?Ͻ=wϽP   P   ��Ͻ�Ͻ�0н�gн�нңн��нێнgн0нE�Ͻh�Ͻ>mϽ�7Ͻ�Ͻ8�νL�ν�Ͻ18Ͻ�mϽP   P   ۜϽ��Ͻ�'нSgн�н=�н(�н�нc�нgн'н�Ͻ�Ͻ�\Ͻ�+ϽnϽVϽ�Ͻq,Ͻ9]ϽP   P   :�Ͻ��Ͻ�н�Tн�н'�нu�н��н�нێнPTн�нt�ϽׁϽ_GϽ0ϽCϽϽeϽiGϽP   P   ;aϽ��Ͻ��Ͻ&0н�pн��нo�нu�н(�н��н�pн�/н��ϽŠϽ�`Ͻ�.Ͻ�ϽϽ�Ͻ�.ϽP   P   �<Ͻ�tϽd�Ͻ\�Ͻ�AнK{н��н'�н=�нңн�zн�Aн��Ͻ��Ͻ�tϽ�<ϽϽ��ν��ν�ϽP   P   3ϽnGϽ�Ͻ)�Ͻ�н�Aн�pн�н�н�н�pн�AнxнL�Ͻ�Ͻ�GϽϽ��ν�νg�νP   P   ��ν�Ͻ�MϽ��Ͻ)�Ͻ\�Ͻ&0н�TнSgн�gн�Tн|0н��Ͻ��Ͻ��Ͻ'NϽ=Ͻ	�ν6�ν�νP   P   R�ν5�ν�Ͻ�MϽ�Ͻd�Ͻ��Ͻ�н�'н�0н(нIн��Ͻ��Ͻ@�Ͻ3NϽϽ��νu�νs�νP   P   �νI�ν5�ν�ϽnGϽ�tϽ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻi�Ͻp�ϽluϽ=HϽ�Ͻ��ν��ν:�νP   P   ��ν`�νe	Ͻ"ϽX4ϽGOϽyjϽL�Ͻ^�ϽP�Ͻ�Ͻ�Ͻm�Ͻ��Ͻ�jϽ�OϽ�4Ͻ�Ͻ�	Ͻ��νP   P   ��ν1�ν�Ͻ�Ͻ&Ͻ�0ϽbDϽ(WϽNgϽ�rϽ�xϽ�xϽsϽ2hϽ�WϽ=EϽ�1ϽϽ[Ͻ�ϽP   P   �	Ͻ�Ͻ�	Ͻ�Ͻ�Ͻ!ϽI,Ͻ�7Ͻ�BϽ�KϽ�PϽRϽ"QϽZLϽ?CϽH8Ͻ�,Ͻ�!ϽiϽ[ϽP   P   �Ͻ�ϽϽ�ϽyϽ� Ͻ$Ͻ�'Ͻ�*Ͻ�-Ͻ&0Ͻ2Ͻ(2Ͻ�0Ͻm.Ͻ�+Ͻ�(Ͻ%Ͻ�!ϽϽP   P   �4Ͻ7Ͻ�7Ͻ�6ϽF4Ͻ�0Ͻ:,Ͻ�'Ͻ�"Ͻ�ϽvϽϽ�Ͻ5ϽϽ�Ͻ�#Ͻ�(Ͻ�,Ͻ�1ϽP   P   �OϽ�WϽ�ZϽ�ZϽ&WϽ-OϽ�DϽ?7Ͻ�*Ͻ�Ͻ�ϽtϽ"	Ͻa	Ͻ�Ͻ+Ͻ�Ͻ�+ϽH8Ͻ=EϽP   P   �jϽzyϽd�ϽA�Ͻ�ϽyϽjϽWϽ�BϽ�-ϽϽrϽϽ%Ͻ5Ͻ�ϽϽm.Ͻ@CϽ�WϽP   P   ��Ͻ �Ͻ,�Ͻ��Ͻ8�ϽЩϽo�Ͻ��ϽBgϽ$KϽ�/Ͻ�Ͻ�Ͻ� Ͻ%Ͻa	Ͻ5Ͻ�0ϽZLϽ2hϽP   P   m�ϽI�Ͻ��Ͻ��ϽF�Ͻ��Ͻ7�Ͻ��Ͻ��Ͻ�rϽ]PϽ�1ϽϽ�ϽϽ"	Ͻ�Ͻ(2Ͻ"QϽsϽP   P   �ϽO�Ͻ�Ͻн�н�нн��Ͻ��Ͻ�Ͻ"xϽ_QϽ�1Ͻ�ϽrϽtϽϽ2ϽRϽ�xϽP   P   �Ͻ,�Ͻ��Ͻн�1нH9н�1н�н��Ͻ��Ͻ�Ͻ"xϽ]PϽ�/ϽϽ�ϽvϽ&0Ͻ�PϽ�xϽP   P   P�Ͻz�Ͻ�нw+н.Hн(Xн�WнHн +н�н��Ͻ�Ͻ�rϽ$KϽ�-Ͻ�Ͻ�Ͻ�-Ͻ�KϽ�rϽP   P   ^�Ͻ��Ͻ��Ͻ+нPн�gн�oн�gн�Oн +н��Ͻ��Ͻ��ϽBgϽ�BϽ�*Ͻ�"Ͻ�*Ͻ�BϽNgϽP   P   L�ϽŴϽ��Ͻ#нAHн�gнxнYxн�gнHн�н��Ͻ��Ͻ��ϽWϽ?7Ͻ�'Ͻ�'Ͻ�7Ͻ(WϽP   P   yjϽh�Ͻ��Ͻ�н�1н�Wн5pнxн�oн�Wн�1нн7�Ͻo�ϽjϽ�DϽ:,Ͻ$ϽI,ϽbDϽP   P   GOϽ�xϽ��ϽA�Ͻ�н�9н�Wн�gн�gн(XнH9н�н��ϽЩϽ
yϽ-OϽ�0Ͻ� Ͻ!Ͻ�0ϽP   P   X4Ͻ�VϽX�Ͻ�Ͻ��Ͻ�н�1нAHнPн.Hн�1н�нF�Ͻ8�Ͻ�Ͻ&WϽF4ϽyϽ�Ͻ&ϽP   P   "Ͻ<6ϽRZϽ��Ͻ�ϽA�Ͻ�н#н+нw+ннн��Ͻ��Ͻ@�Ͻ�ZϽ�6Ͻ�Ͻ�Ͻ�ϽP   P   e	Ͻ2Ͻ�7ϽRZϽX�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�н��Ͻ�Ͻ��Ͻ,�Ͻd�Ͻ�ZϽ�7ϽϽ�	Ͻ�ϽP   P   `�ν�Ͻ2Ͻ<6Ͻ�VϽ�xϽh�ϽŴϽ��Ͻz�Ͻ,�ϽO�ϽI�Ͻ �ϽzyϽ�WϽ7Ͻ�Ͻ�Ͻ1�νP   P   �Ͻ� ϽW)Ͻ�7Ͻ[IϽI\Ͻ�oϽ�Ͻ�Ͻ�Ͻt�ϽR�Ͻ�Ͻo�Ͻ1pϽ�\Ͻ�IϽ�7Ͻ�)Ͻ� ϽP   P   � Ͻ� Ͻ�$Ͻ,-Ͻ�8Ͻ�FϽ�TϽcϽ�nϽTwϽ\|ϽA|Ͻ�wϽoϽ�cϽ�UϽ<GϽT9Ͻ�-Ͻ�$ϽP   P   �)Ͻ�(Ͻ�)Ͻ	-Ͻ�2Ͻ�:ϽFCϽ�KϽdSϽ�XϽ^Ͻ�_ϽC^ϽKYϽ�SϽLϽ�CϽ;ϽE3Ͻ�-ϽP   P   �7Ͻr6ϽG6Ͻ�7Ͻ�8Ͻ�:Ͻ�<Ͻ}?ϽqBϽ�DϽ{FϽ!GϽXGϽ�FϽ*EϽ#CϽ4@Ͻ�=Ͻ;ϽT9ϽP   P   �IϽhKϽ�JϽGKϽrIϽrFϽ9CϽ�?Ͻu<Ͻ�9ϽO7Ͻ5Ͻ�4Ͻ�5Ͻ�7Ͻ*:Ͻ�<Ͻ4@Ͻ�CϽ<GϽP   P   �\Ͻ�bϽ�eϽ�eϽ`bϽ3\Ͻ�TϽ�KϽZBϽw9Ͻl1Ͻ ,Ͻ�)Ͻ�)ϽJ,Ͻ�1Ͻ*:Ͻ#CϽLϽ�UϽP   P   1pϽ�{Ͻ��Ͻ�Ͻx�ϽR{Ͻ�oϽ�bϽfSϽ�DϽ\7Ͻ�+Ͻ�$Ͻ^#Ͻ=%ϽJ,Ͻ�7Ͻ+EϽ�SϽ�cϽP   P   o�Ͻv�ϽC�Ͻ��ϽQ�Ͻ��Ͻ��ϽׁϽ�nϽbXϽ%FϽ35Ͻ�)Ͻ^#Ͻ^#Ͻ�)Ͻ�5Ͻ�FϽKYϽoϽP   P   �Ͻ��Ͻ@�Ͻ��Ͻ#�Ͻ��Ͻ�Ͻ4�Ͻ��Ͻ�vϽ�]Ͻ�FϽF4Ͻ�)Ͻ�$Ͻ�)Ͻ�4ϽXGϽD^Ͻ�wϽP   P   R�Ͻ��ϽB�Ͻz�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�ϽՙϽ�{Ͻ#_Ͻ�FϽ35Ͻ�+Ͻ ,Ͻ5Ͻ!GϽ�_ϽA|ϽP   P   t�Ͻ|�Ͻ_�ϽE�Ͻ�нAн�н�Ͻ�Ͻ�Ͻ؜Ͻ�{Ͻ�]Ͻ%FϽ\7Ͻl1ϽO7Ͻ{FϽ^Ͻ\|ϽP   P   �Ͻt�Ͻ!�ϽF�ϽRн�н�нн��Ͻ��Ͻ�ϽՙϽ�vϽbXϽ�DϽw9Ͻ�9Ͻ�DϽ�XϽTwϽP   P   �Ͻx�Ͻa�Ͻ%�Ͻ�н+нm1нq+н�н��Ͻ�Ͻ�Ͻ��Ͻ�nϽfSϽZBϽu<ϽqBϽdSϽ�nϽP   P   �ϽG�Ͻ��Ͻ<�Ͻ?н�+нU7нc7нq+нн�Ͻ��Ͻ4�ϽׁϽ�bϽ�KϽ�?Ͻ}?Ͻ�KϽcϽP   P   �oϽ�Ͻ6�Ͻ=�Ͻ�н�нl1нU7нm1н�н�н�Ͻ�Ͻ��Ͻ�oϽ�TϽ9CϽ�<ϽFCϽ�TϽP   P   I\Ͻ&{Ͻ�Ͻ��Ͻ��ϽEн�н�+н+н�нAн��Ͻ��Ͻ��ϽR{Ͻ3\ϽrFϽ�:Ͻ�:Ͻ�FϽP   P   [IϽNbϽq�Ͻ:�Ͻ0�Ͻ��Ͻ�н?н�нRн�н��Ͻ#�ϽQ�Ͻx�Ͻ`bϽrIϽ�8Ͻ�2Ͻ�8ϽP   P   �7Ͻ�JϽ�eϽǅϽ:�Ͻ��Ͻ=�Ͻ<�Ͻ%�ϽF�ϽE�Ͻz�Ͻ��Ͻ��Ͻ�Ͻ�eϽFKϽ�7Ͻ	-Ͻ,-ϽP   P   W)Ͻ6Ͻ�JϽ�eϽq�Ͻ�Ͻ6�Ͻ��Ͻ`�Ͻ!�Ͻ_�ϽB�Ͻ@�ϽC�Ͻ��Ͻ�eϽ�JϽG6Ͻ�)Ͻ�$ϽP   P   � Ͻ�(Ͻ6Ͻ�JϽNbϽ&{Ͻ�ϽG�Ͻx�Ͻt�Ͻ|�Ͻ��Ͻ��Ͻv�Ͻ�{Ͻ�bϽhKϽr6Ͻ�(Ͻ� ϽP   P   78Ͻ�:Ͻ^AϽ�KϽ8XϽ�gϽvϽ�Ͻ��ϽH�ϽϖϽL�Ͻ�Ͻ��ϽPvϽ�gϽ�XϽ�KϽ�AϽ�:ϽP   P   �:Ͻ�:Ͻ>Ͻ�DϽ}LϽ�VϽ�aϽ�kϽ�tϽ�zϽ)~Ͻ~ϽL{Ͻ�tϽ�kϽ.bϽ2WϽ�LϽ�DϽQ>ϽP   P   �AϽ�@Ͻ�AϽ_DϽ�HϽNϽ{TϽ	[ϽS`Ͻ@eϽ�gϽ�hϽhϽ�eϽ�`Ͻ}[Ͻ�TϽ�NϽIϽ�DϽP   P   �KϽ"KϽ�JϽ�KϽ�LϽ@NϽPϽRϽ�SϽ�UϽ�VϽ9WϽ_WϽ�VϽ�UϽ�SϽ�RϽ�PϽ�NϽ�LϽP   P   �XϽvZϽl[ϽVZϽ�XϽ�VϽ�TϽ�QϽ�NϽ�LϽ�JϽJϽ�IϽ?JϽNKϽ MϽ�OϽ�RϽ�TϽ2WϽP   P   �gϽgkϽ�mϽ�mϽ�jϽ{gϽ�aϽ�ZϽ�SϽfLϽ^GϽ�CϽ�AϽ�AϽDϽ�GϽ MϽ�SϽ}[Ͻ.bϽP   P   PvϽϽJ�Ͻ��Ͻ<�Ͻ�~ϽvϽLkϽr`Ͻ@UϽ'KϽ�CϽ>Ͻ%<Ͻb>ϽDϽNKϽ�UϽ�`Ͻ�kϽP   P   ��Ͻ-�Ͻ<�Ͻ\�ϽC�Ͻ�Ͻ��Ͻ�ϽNtϽeϽ�VϽ�IϽ�AϽ<<Ͻ%<Ͻ�AϽ?JϽ�VϽ�eϽ�tϽP   P   �ϽݞϽ�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ{zϽ�gϽ�VϽ�IϽ�AϽ>Ͻ�AϽ�IϽ_WϽhϽL{ϽP   P   L�Ͻ��Ͻ��Ͻs�Ͻ��Ͻ��ϽS�Ͻ	�Ͻ*�Ͻ�Ͻ�}ϽYhϽ�VϽ�IϽ�CϽ�CϽJϽ9WϽ�hϽ~ϽP   P   ϖϽw�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽҮϽ��Ͻ�}Ͻ�gϽ�VϽ'KϽ^GϽ�JϽ�VϽ�gϽ)~ϽP   P   H�Ͻ�Ͻ�Ͻ%�Ͻ��Ͻ��Ͻ��Ͻx�Ͻ��Ͻ��ϽҮϽ�Ͻ{zϽeϽ@UϽfLϽ�LϽ�UϽ@eϽ�zϽP   P   ��Ͻ��Ͻ��ϽK�Ͻ�Ͻ^�ϽRнN�Ͻ)�Ͻ��Ͻ��Ͻ*�Ͻ��ϽNtϽr`Ͻ�SϽ�NϽ�SϽS`Ͻ�tϽP   P   �ϽȞϽ[�Ͻ��Ͻ��Ͻp�Ͻr	н	нN�Ͻx�Ͻ��Ͻ	�Ͻ��Ͻ�ϽLkϽ�ZϽ�QϽRϽ	[Ͻ�kϽP   P   vϽ�Ͻ��Ͻ~�Ͻ��Ͻ��Ͻнr	нRн��Ͻ��ϽS�Ͻ�Ͻ��ϽvϽ�aϽ�TϽPϽ{TϽ�aϽP   P   �gϽ�~Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻp�Ͻ^�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�~Ͻ{gϽ�VϽ@NϽNϽ�VϽP   P   8XϽkϽ��ϽF�Ͻ0�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��ϽC�Ͻ<�Ͻ�jϽ�XϽ�LϽ�HϽ}LϽP   P   �KϽ]ZϽ�mϽ��ϽF�Ͻ��Ͻ~�Ͻ��ϽK�Ͻ%�Ͻ��Ͻs�Ͻ�Ͻ\�Ͻ��Ͻ�mϽVZϽ�KϽ_DϽ�DϽP   P   ^AϽ�JϽ�ZϽ�mϽ��Ͻ�Ͻ��Ͻ[�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ<�ϽJ�Ͻ�mϽl[Ͻ�JϽ�AϽ>ϽP   P   �:Ͻ�@Ͻ�JϽ]ZϽkϽ�~Ͻ�ϽȞϽ��Ͻ�Ͻw�Ͻ��ϽݞϽ-�ϽϽgkϽvZϽ"KϽ�@Ͻ�:ϽP   P   �MϽ�NϽ�SϽ [Ͻ�dϽpϽSzϽV�Ͻ_�Ͻ��Ͻ��Ͻ��Ͻ݋ϽфϽ�zϽ:pϽ�eϽh[Ͻ�SϽ�NϽP   P   �NϽ�NϽ$QϽ�UϽ`\Ͻ�cϽ3kϽ�rϽsyϽ(~Ͻ��Ͻ׀Ͻj~ϽTyϽ	sϽ�kϽdϽ|\Ͻ�UϽCQϽP   P   �SϽSϽ�SϽsUϽYϽ*]ϽeaϽgfϽ�jϽ�nϽFpϽ_qϽfpϽ�nϽgkϽ�fϽ bϽ�]Ͻ�YϽ�UϽP   P   h[Ͻl[ϽT[ϽG[Ͻ[\Ͻe]Ͻm^Ͻ�_ϽaϽ�bϽ;cϽodϽodϽxcϽ�bϽ<aϽ(`Ͻ�^Ͻ�]Ͻ|\ϽP   P   �eϽ�eϽLfϽ�eϽVeϽ�cϽtaϽ�_Ͻp^Ͻ]Ͻ�ZϽEZϽsZϽ�ZϽ�ZϽ9]Ͻ&_Ͻ(`Ͻ bϽdϽP   P   :pϽ&sϽ[tϽBtϽ�rϽpϽMkϽDfϽ?aϽ�\Ͻ�XϽDUϽ&SϽ6SϽMUϽYϽ9]Ͻ<aϽ�fϽ�kϽP   P   �zϽ�Ͻ��Ͻq�Ͻ��Ͻ�ϽXzϽ�rϽ�jϽ0bϽ�ZϽ#UϽUQϽ�PϽ�QϽMUϽ�ZϽ�bϽgkϽ	sϽP   P   фϽ��Ͻ��Ͻ��ϽȗϽǓϽ��Ͻd�Ͻ7yϽ�nϽ cϽ(ZϽ�RϽ�PϽ�PϽ6SϽ�ZϽxcϽ�nϽTyϽP   P   ݋Ͻ��Ͻ��Ͻ/�Ͻ�Ͻ�Ͻ\�Ͻ��Ͻa�Ͻ�}ϽpϽdϽjZϽ�RϽUQϽ&SϽsZϽodϽfpϽj~ϽP   P   ��Ͻ��ϽB�Ͻ�Ͻ!�Ͻ�Ͻ�Ͻ��ϽV�Ͻ��Ͻg�ϽqϽdϽ(ZϽ#UϽDUϽEZϽodϽ_qϽ׀ϽP   P   ��Ͻ�Ͻ>�Ͻ�Ͻ\�Ͻ)�Ͻ!�Ͻ�Ͻ0�Ͻ��Ͻq�Ͻg�ϽpϽ cϽ�ZϽ�XϽ�ZϽ;cϽFpϽ��ϽP   P   ��ϽӤϽ �Ͻq�Ͻ��Ͻz�Ͻ��Ͻ(�Ͻ@�Ͻ�Ͻ��Ͻ��Ͻ�}Ͻ�nϽ0bϽ�\Ͻ]Ͻ�bϽ�nϽ(~ϽP   P   _�Ͻ��Ͻ-�Ͻ��Ͻ$�Ͻ��Ͻ��Ͻ�ϽJ�Ͻ@�Ͻ0�ϽV�Ͻa�Ͻ7yϽ�jϽ?aϽp^ϽaϽ�jϽsyϽP   P   V�ϽŘϽ�Ͻ.�ϽL�Ͻ�Ͻ��Ͻd�Ͻ�Ͻ(�Ͻ�Ͻ��Ͻ��Ͻd�Ͻ�rϽDfϽ�_Ͻ�_ϽgfϽ�rϽP   P   SzϽ��Ͻ	�Ͻ3�Ͻ�Ͻ��Ͻ!�Ͻ��Ͻ��Ͻ��Ͻ!�Ͻ�Ͻ\�Ͻ��ϽXzϽMkϽtaϽm^ϽeaϽ3kϽP   P   pϽ�ϽؓϽ!�Ͻ/�Ͻ	�Ͻ��Ͻ�Ͻ��Ͻz�Ͻ)�Ͻ�Ͻ�ϽǓϽ�ϽpϽ�cϽe]Ͻ*]Ͻ�cϽP   P   �dϽ�rϽS�ϽėϽ��Ͻ/�Ͻ�ϽL�Ͻ$�Ͻ��Ͻ\�Ͻ!�Ͻ�ϽȗϽ��Ͻ�rϽVeϽ[\ϽYϽ`\ϽP   P    [Ͻ�eϽDtϽR�ϽėϽ!�Ͻ3�Ͻ.�Ͻ��Ͻq�Ͻ�Ͻ�Ͻ/�Ͻ��Ͻq�ϽBtϽ�eϽG[ϽsUϽ�UϽP   P   �SϽI[Ͻ�eϽDtϽS�ϽؓϽ	�Ͻ�Ͻ-�Ͻ �Ͻ>�ϽB�Ͻ��Ͻ��Ͻ��Ͻ[tϽLfϽT[Ͻ�SϽ$QϽP   P   �NϽ�RϽI[Ͻ�eϽ�rϽ�Ͻ��ϽŘϽ��ϽӤϽ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ&sϽ�eϽl[ϽSϽ�NϽP   P   �\Ͻ ^Ͻ�aϽkgϽnϽ�uϽc~Ͻ��ϽY�Ͻ~�Ͻ�Ͻa�Ͻ��ϽӅϽ�~Ͻ&vϽ�nϽ�gϽ�aϽ^ϽP   P   ^Ͻ�]Ͻ>`Ͻ.cϽhϽ@mϽsϽ�xϽA}Ͻ3�Ͻ�Ͻ0�Ͻ7�Ͻg}Ͻ�xϽNsϽEmϽ�gϽtcϽ=`ϽP   P   �aϽ�`Ͻ�aϽUcϽ`eϽ�hϽLlϽpϽ�rϽ�tϽ�vϽ�wϽ�vϽ�tϽ(sϽIpϽ�lϽ�hϽ�eϽtcϽP   P   �gϽgϽ gϽcgϽ�gϽ�hϽ	jϽ�jϽwkϽ�lϽ&mϽmϽ�lϽ�mϽ�lϽ�kϽ�jϽ�iϽ�hϽ�gϽP   P   �nϽoϽ�nϽ�nϽOnϽ-mϽ\lϽ�jϽ�hϽ�gϽ�gϽgϽ�eϽ gϽ�gϽ�gϽ�iϽ�jϽ�lϽFmϽP   P   &vϽ�xϽmzϽFzϽ�xϽ�uϽ/sϽpϽ�kϽ�gϽ6dϽ�bϽ�aϽ�aϽ�bϽ�dϽ�gϽ�kϽIpϽNsϽP   P   �~Ͻ��Ͻ��Ͻ؆Ͻ��Ͻ��ϽF~Ͻ�xϽ[rϽ[lϽmgϽ�bϽ`Ͻ�^ϽF`Ͻ�bϽ�gϽ�lϽ(sϽ�xϽP   P   ӅϽ}�ϽD�Ͻ��Ͻ��Ͻ�Ͻ�Ͻm�Ͻ7}Ͻ�tϽ1mϽ�fϽ�aϽ�^Ͻ�^Ͻ�aϽ gϽ�mϽ�tϽg}ϽP   P   ��Ͻ"�ϽA�Ͻ}�Ͻ[�Ͻ��ϽכϽ�Ͻ�Ͻ��ϽvϽ�lϽ�eϽ�aϽ`Ͻ�aϽ�eϽ�lϽ�vϽ7�ϽP   P   a�ϽT�Ͻ-�Ͻ��ϽP�Ͻ�Ͻ��ϽݣϽ)�ϽE�Ͻ��Ͻ�wϽ�lϽ�fϽ�bϽ�bϽgϽmϽ�wϽ0�ϽP   P   �Ͻ˝ϽI�Ͻ1�Ͻ��ϽR�Ͻt�ϽB�Ͻ��Ͻ��Ͻ��Ͻ��ϽvϽ1mϽmgϽ6dϽ�gϽ&mϽ�vϽ�ϽP   P   ~�ϽɝϽ��Ͻt�Ͻ��Ͻ��Ͻ�Ͻ��ϽH�Ͻ��Ͻ��ϽE�Ͻ��Ͻ�tϽ[lϽ�gϽ�gϽ�lϽ�tϽ3�ϽP   P   Y�Ͻ �Ͻ5�Ͻ[�Ͻ��ϽF�Ͻ��ϽH�Ͻ��ϽH�Ͻ��Ͻ)�Ͻ�Ͻ7}Ͻ[rϽ�kϽ�hϽwkϽ�rϽA}ϽP   P   ��ϽG�Ͻ��ϽJ�Ͻ¿Ͻ��Ͻw�ϽB�ϽH�Ͻ��ϽB�ϽݣϽ�Ͻm�Ͻ�xϽpϽ�jϽ�jϽpϽ�xϽP   P   c~Ͻs�Ͻ�Ͻ��Ͻl�Ͻ�Ͻs�Ͻw�Ͻ��Ͻ�Ͻt�Ͻ��ϽכϽ�ϽF~Ͻ/sϽ\lϽ	jϽLlϽsϽP   P   �uϽ��Ͻ�Ͻ��Ͻ4�Ͻ\�Ͻ�Ͻ��ϽF�Ͻ��ϽR�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ�uϽ-mϽ�hϽ�hϽ@mϽP   P   nϽ�xϽ��Ͻ��Ͻ.�Ͻ4�Ͻl�Ͻ¿Ͻ��Ͻ��Ͻ��ϽP�Ͻ[�Ͻ��Ͻ��Ͻ�xϽOnϽ�gϽ`eϽhϽP   P   kgϽoϽBzϽ��Ͻ��Ͻ��Ͻ��ϽJ�Ͻ[�Ͻt�Ͻ1�Ͻ��Ͻ}�Ͻ��Ͻ؆ϽFzϽ�nϽbgϽUcϽ.cϽP   P   �aϽgϽ�nϽBzϽ��Ͻ�Ͻ�Ͻ��Ͻ5�Ͻ��ϽI�Ͻ-�ϽA�ϽD�Ͻ��ϽmzϽ�nϽ gϽ�aϽ>`ϽP   P    ^Ͻ�`ϽgϽoϽ�xϽ��Ͻs�ϽG�Ͻ �ϽɝϽ˝ϽT�Ͻ"�Ͻ}�Ͻ��Ͻ�xϽoϽgϽ�`Ͻ�]ϽP   P   �hϽ-jϽ�lϽ�pϽ�uϽ'|ϽˁϽ͆Ͻw�Ͻ��Ͻ��Ͻ��Ͻ��ϽˆϽ�Ͻo|Ͻ%vϽ�pϽ�lϽ6jϽP   P   6jϽ#jϽkϽ�mϽGqϽxuϽ�yϽm}Ͻ[�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻw}Ͻ�yϽ�uϽgqϽ�mϽkϽP   P   �lϽ�lϽilϽ�mϽ�oϽ�qϽ&tϽwvϽOyϽb{Ͻ�|Ͻ�|Ͻ�|Ͻ\{Ͻ�yϽ�vϽ�tϽrϽ�oϽ�mϽP   P   �pϽ�pϽ�pϽ�pϽ5qϽ�qϽbrϽ&sϽFtϽ�tϽZuϽ�uϽ�uϽ�uϽ�tϽqtϽNsϽjrϽrϽgqϽP   P   %vϽ�vϽ(wϽ�vϽ�uϽ�uϽtϽsϽwrϽ`qϽ�pϽ�oϽ)pϽ�oϽ�pϽ�qϽ�rϽNsϽ�tϽ�uϽP   P   o|ϽS}Ͻ2~Ͻ"~ϽU}Ͻ'|Ͻ�yϽvvϽFtϽ`qϽGoϽHmϽ�lϽ�lϽWmϽtoϽ�qϽqtϽ�vϽ�yϽP   P   �Ͻz�Ͻ��ϽH�Ͻ|�Ͻs�Ͻ��Ͻp}ϽyϽ�tϽ~pϽBmϽ�kϽPjϽ�kϽWmϽ�pϽ�tϽ�yϽw}ϽP   P   ˆϽa�Ͻ)�Ͻ��Ͻ��Ͻ�ϽY�Ͻ��Ͻv�ϽE{ϽzuϽ�oϽ�lϽEjϽPjϽ�lϽ�oϽ�uϽ\{Ͻ��ϽP   P   ��Ͻ��Ͻ^�ϽP�Ͻ*�Ͻo�Ͻ�Ͻ��Ͻ2�Ͻ��ϽL|Ͻ�uϽ�oϽ�lϽ�kϽ�lϽ)pϽ�uϽ�|Ͻ��ϽP   P   ��Ͻ��Ͻ՝Ͻ��Ͻ��Ͻ[�Ͻm�ϽʝϽ��Ͻy�Ͻ��Ͻ�|Ͻ�uϽ�oϽBmϽHmϽ�oϽ�uϽ�|Ͻ��ϽP   P   ��Ͻt�Ͻ��Ͻ`�Ͻ�Ͻ�Ͻ�Ͻ_�Ͻ=�Ͻa�Ͻ;�Ͻ��ϽL|ϽzuϽ~pϽGoϽ�pϽZuϽ�|Ͻ��ϽP   P   ��Ͻ~�Ͻ�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ�ϽԫϽ�Ͻa�Ͻy�Ͻ��ϽE{Ͻ�tϽ`qϽ`qϽ�tϽb{Ͻ��ϽP   P   w�Ͻ��Ͻ��Ͻ۫Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽԫϽ=�Ͻ��Ͻ2�Ͻv�ϽyϽFtϽwrϽFtϽOyϽ[�ϽP   P   ͆Ͻ֑ϽĝϽf�Ͻ�Ͻ��ϽN�Ͻo�Ͻ��Ͻ�Ͻ_�ϽʝϽ��Ͻ��Ͻp}ϽvvϽsϽ&sϽwvϽm}ϽP   P   ˁϽ �Ͻk�Ͻj�Ͻ3�Ͻi�Ͻ#�ϽN�Ͻ�Ͻ��Ͻ�Ͻm�Ͻ�ϽY�Ͻ��Ͻ�yϽtϽbrϽ&tϽ�yϽP   P   '|Ͻ��Ͻ�Ͻ<�Ͻf�Ͻ �Ͻi�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ[�Ͻo�Ͻ�Ͻs�Ͻ'|Ͻ�uϽ�qϽ�qϽxuϽP   P   �uϽ:}Ͻ|�Ͻ��ϽC�Ͻf�Ͻ3�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ*�Ͻ��Ͻ|�ϽU}Ͻ�uϽ5qϽ�oϽGqϽP   P   �pϽ�vϽ~ϽH�Ͻ��Ͻ<�Ͻj�Ͻf�Ͻ۫Ͻ�Ͻ`�Ͻ��ϽP�Ͻ��ϽH�Ͻ"~Ͻ�vϽ�pϽ�mϽ�mϽP   P   �lϽ�pϽwϽ~Ͻ|�Ͻ�Ͻk�ϽĝϽ��Ͻ�Ͻ��Ͻ՝Ͻ^�Ͻ)�Ͻ��Ͻ2~Ͻ(wϽ�pϽilϽkϽP   P   -jϽHlϽ�pϽ�vϽ9}Ͻ��Ͻ �Ͻ֑Ͻ��Ͻ~�Ͻt�Ͻ��Ͻ��Ͻa�Ͻz�ϽS}Ͻ�vϽ�pϽ�lϽ#jϽP   P   RrϽ#sϽKuϽ)xϽD|Ͻ)�Ͻ7�Ͻ�Ͻ��Ͻ��Ͻ�ϽԍϽ��ϽĈϽV�Ͻ��Ͻ�{Ͻ?xϽ9uϽ2sϽP   P   2sϽOsϽ�sϽ�uϽbxϽm{Ͻ�~Ͻ��Ͻ8�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ��ϽE�Ͻ Ͻ�{Ͻ�xϽ"vϽ,tϽP   P   9uϽ�tϽuϽ
vϽewϽyϽ�zϽ}|ϽV~Ͻ�Ͻ��Ͻ$�Ͻ��Ͻ�ϽF~Ͻ�|Ͻ�zϽ5yϽ#wϽ"vϽP   P   ?xϽ�wϽ�wϽJxϽExϽ yϽ�yϽ"zϽ�zϽ�zϽ{Ͻ�{Ͻ�{Ͻ{Ͻ�zϽ�zϽvzϽ�yϽ5yϽ�xϽP   P   �{Ͻ�|Ͻb|Ͻ~|Ͻ|Ͻ�{Ͻ�zϽ1zϽpyϽRxϽ"xϽ�wϽ0xϽ�wϽ-xϽ�xϽMyϽvzϽ�zϽ�{ϽP   P   ��Ͻ�Ͻ��Ͻ��Ͻ��ϽY�Ͻ�~Ͻ�|Ͻ�zϽnxϽ�wϽ�uϽ�tϽ�tϽ�uϽ�wϽ�xϽ�zϽ�|Ͻ ϽP   P   V�Ͻ��ϽшϽ��Ͻ�Ͻ��ϽJ�Ͻ�ϽR~Ͻ�zϽxϽ�uϽntϽLtϽ8tϽ�uϽ-xϽ�zϽF~ϽE�ϽP   P   ĈϽ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ1�ϽgϽ{Ͻ]wϽ�tϽ�sϽLtϽ�tϽ�wϽ{Ͻ�Ͻ��ϽP   P   ��Ͻ)�Ͻ��Ͻ��Ͻ)�Ͻ��Ͻ��ϽƐϽ��Ͻ�Ͻl�Ͻ�{Ͻ,xϽ�tϽntϽ�tϽ0xϽ�{Ͻ��Ͻ�ϽP   P   ԍϽ�Ͻq�ϽϝϽq�Ͻ`�Ͻ}�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ�{Ͻ]wϽ�uϽ�uϽ�wϽ�{Ͻ$�Ͻ��ϽP   P   �ϽٕϽe�Ͻ��Ͻh�ϽM�Ͻ��Ͻ_�ϽP�Ͻ��ϽɏϽ��Ͻl�Ͻ{ϽxϽ�wϽ"xϽ{Ͻ��Ͻ�ϽP   P   ��Ͻ��Ͻ�ϽL�Ͻ]�ϽM�Ͻ�Ͻg�ϽB�Ͻ؜Ͻ��Ͻ��Ͻ�ϽgϽ�zϽnxϽRxϽ�zϽ�Ͻ�ϽP   P   ��Ͻ#�Ͻj�ϽS�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ|�ϽB�ϽP�Ͻ�Ͻ��Ͻ1�ϽR~Ͻ�zϽpyϽ�zϽV~Ͻ8�ϽP   P   �Ͻ��Ͻ}�ϽL�Ͻw�Ͻz�Ͻ�ϽO�Ͻ��Ͻg�Ͻ_�Ͻ��ϽƐϽ��Ͻ�Ͻ�|Ͻ1zϽ"zϽ}|Ͻ��ϽP   P   7�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ}�Ͻ��Ͻ��ϽJ�Ͻ�~Ͻ�zϽ�yϽ�zϽ�~ϽP   P   )�Ͻ��Ͻ�Ͻx�ϽT�ϽP�Ͻ�Ͻz�Ͻ��ϽM�ϽM�Ͻ`�Ͻ��Ͻ�Ͻ��ϽY�Ͻ�{Ͻ yϽyϽm{ϽP   P   D|ϽŁϽϽ��Ͻx�ϽT�Ͻ��Ͻw�Ͻ��Ͻ]�Ͻh�Ͻq�Ͻ)�Ͻ��Ͻ�Ͻ��Ͻ|ϽExϽewϽbxϽP   P   )xϽY|Ͻq�Ͻ�Ͻ��Ͻx�Ͻ��ϽL�ϽS�ϽL�Ͻ��ϽϝϽ��Ͻ�Ͻ��Ͻ��Ͻ~|ϽJxϽ
vϽ�uϽP   P   KuϽ�wϽ�|Ͻq�ϽϽ�Ͻ�Ͻ}�Ͻj�Ͻ�Ͻe�Ͻq�Ͻ��Ͻ�ϽшϽ��Ͻb|Ͻ�wϽuϽ�sϽP   P   #sϽ�tϽ�wϽY|ϽŁϽ��Ͻ��Ͻ��Ͻ#�Ͻ��ϽٕϽ�Ͻ)�Ͻ��Ͻ��Ͻ�Ͻ�|Ͻ�wϽ�tϽOsϽP   P   czϽszϽU|Ͻh~Ͻ\�Ͻ'�Ͻ�Ͻ��ϽیϽ�Ͻv�Ͻ�Ͻ��Ͻ��ϽЇϽq�Ͻ �Ͻ~Ͻ,|ϽqzϽP   P   qzϽ�zϽu{Ͻ�|Ͻ�~Ͻm�ϽN�ϽP�Ͻ׆Ͻ�Ͻ8�Ͻ�Ͻ*�Ͻ�Ͻ��ϽB�Ͻ��ϽϽ�|Ͻ�{ϽP   P   ,|Ͻ�{ϽG|Ͻ�|Ͻ�}Ͻ�~Ͻa�Ͻ��Ͻ��Ͻ-�Ͻ��Ͻ�ϽǄϽ=�Ͻ��Ͻ��Ͻ7�Ͻ�~ϽR}Ͻ�|ϽP   P   ~Ͻ�~Ͻn~Ͻ�~Ͻ�~Ͻ�~Ͻ#ϽgϽL�Ͻ��Ͻ��Ͻ��Ͻ܀Ͻ�Ͻ�ϽZ�Ͻ�Ͻ_Ͻ�~ϽϽP   P    �ϽS�Ͻs�ϽG�Ͻ7�Ͻ��ϽW�Ͻ�Ͻ�~ϽZ~Ͻ�~Ͻ�~Ͻ�}Ͻ�~Ͻ�~Ͻ�~Ͻ�~Ͻ�Ͻ7�Ͻ��ϽP   P   q�ϽԅϽ��Ͻ��Ͻ_�Ͻ[�Ͻ�ϽϽ�Ͻj~Ͻ�|ϽI|Ͻ|Ͻ�{Ͻ�|Ͻ{|Ͻ�~ϽZ�Ͻ��ϽB�ϽP   P   ЇϽ��Ͻ9�ϽS�Ͻ\�Ͻ��Ͻ��ϽY�Ͻ��ϽހϽ�~Ͻ~|Ͻp{Ͻ�zϽ{Ͻ�|Ͻ�~Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ�Ͻ=�Ͻ��Ͻ_�Ͻ-�Ͻ��Ͻ��ϽÆϽ�Ͻ߀Ͻ�~Ͻ|Ͻ_zϽ�zϽ�{Ͻ�~Ͻ�Ͻ=�Ͻ�ϽP   P   ��Ͻ͐Ͻ-�Ͻ.�Ͻ,�Ͻ%�Ͻ\�Ͻh�Ͻ�Ͻ�ϽބϽ��Ͻ�}Ͻ|Ͻp{Ͻ|Ͻ�}Ͻ܀ϽǄϽ*�ϽP   P   �Ͻ��ϽÕϽ��Ͻ&�ϽI�ϽM�Ͻ�Ͻs�Ͻ؍Ͻ�Ͻ��Ͻ��Ͻ�~Ͻ~|ϽI|Ͻ�~Ͻ��Ͻ�Ͻ�ϽP   P   v�ϽޓϽ�Ͻ��Ͻ�Ͻ�Ͻ,�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�ϽބϽ߀Ͻ�~Ͻ�|Ͻ�~Ͻ��Ͻ��Ͻ8�ϽP   P   �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽJ�ϽءϽ��Ͻ˙Ͻ��Ͻ؍Ͻ�Ͻ�ϽހϽj~ϽZ~Ͻ��Ͻ-�Ͻ�ϽP   P   یϽ��Ͻ�Ͻ��ϽâϽZ�Ͻ��Ͻ6�Ͻ��Ͻ��Ͻ�Ͻs�Ͻ�ϽÆϽ��Ͻ�Ͻ�~ϽL�Ͻ��Ͻ׆ϽP   P   ��ϽT�Ͻ�Ͻ��ϽǡϽ�Ͻe�Ͻ��Ͻ6�ϽءϽ��Ͻ�Ͻh�Ͻ��ϽY�ϽϽ�ϽgϽ��ϽP�ϽP   P   �ϽϽ^�Ͻt�Ͻ9�ϽX�Ͻb�Ͻe�Ͻ��ϽJ�Ͻ,�ϽM�Ͻ\�Ͻ��Ͻ��Ͻ�ϽW�Ͻ#Ͻa�ϽN�ϽP   P   '�Ͻ��Ͻ1�Ͻ �Ͻ�Ͻ�ϽX�Ͻ�ϽZ�Ͻ��Ͻ�ϽI�Ͻ%�Ͻ-�Ͻ��Ͻ[�Ͻ��Ͻ�~Ͻ�~Ͻm�ϽP   P   \�Ͻ��ϽM�Ͻi�ϽY�Ͻ�Ͻ9�ϽǡϽâϽ��Ͻ�Ͻ&�Ͻ,�Ͻ_�Ͻ\�Ͻ_�Ͻ7�Ͻ�~Ͻ�}Ͻ�~ϽP   P   h~Ͻ�Ͻs�Ͻ`�Ͻi�Ͻ �Ͻt�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ.�Ͻ��ϽS�Ͻ��ϽG�Ͻ�~Ͻ�|Ͻ�|ϽP   P   U|Ͻm~Ͻ��Ͻs�ϽM�Ͻ1�Ͻ^�Ͻ�Ͻ�Ͻ��Ͻ�ϽÕϽ-�Ͻ=�Ͻ9�Ͻ��Ͻs�Ͻn~ϽG|Ͻu{ϽP   P   szϽ�{Ͻm~Ͻ�Ͻ��Ͻ��ϽϽT�Ͻ��Ͻ��ϽޓϽ��Ͻ͐Ͻ�Ͻ��ϽԅϽS�Ͻ�~Ͻ�{Ͻ�zϽP   P   i�Ͻ��Ͻt�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��ϽӍϽ��Ͻ�ϽƇϽ}�Ͻ�ϽS�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ́Ͻ��Ͻ1�Ͻ��Ͻ-�Ͻ�ϽʊϽS�Ͻx�ϽȊϽ�Ͻw�Ͻ��Ͻf�Ͻ��Ͻ�Ͻ5�ϽP   P   S�Ͻo�Ͻ~�ϽفϽ��Ͻ݃Ͻ�Ͻ��ϽφϽk�Ͻ��Ͻ�Ͻ��Ͻz�Ͻ��Ͻ��Ͻ�ϽރϽ��Ͻ�ϽP   P   �ϽK�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ̃Ͻ`�Ͻo�Ͻo�Ͻz�Ͻ5�Ͻ<�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽރϽ��ϽP   P   }�Ͻ��Ͻ�Ͻ��Ͻ��ϽN�ϽфϽ��Ͻ\�Ͻ�Ͻ��ϽقϽz�Ͻ�ϽςϽ5�Ͻ<�Ͻ��Ͻ�Ͻf�ϽP   P   ƇϽK�Ͻ�Ͻ�Ͻ,�Ͻ��Ͻ��Ͻ��ϽF�Ͻ�Ͻ��ϽϽ�ϽՁϽ�Ͻ҂Ͻ5�Ͻ��Ͻ��Ͻ��ϽP   P   �Ͻ4�Ͻ'�ϽȌϽ'�Ͻ6�ϽމϽE�ϽϽ��Ͻ؂Ͻ�Ͻx�Ͻ�Ͻl�Ͻ�ϽςϽ��Ͻ��Ͻw�ϽP   P   ��Ͻ֍Ͻ��Ͻs�Ͻw�Ͻ��Ͻ��Ͻ��Ͻ�ϽG�Ͻj�ϽׂϽ߁Ͻ׀Ͻ�ϽՁϽ�Ͻ��Ͻz�Ͻ�ϽP   P   ӍϽ��Ͻ�ϽM�Ͻ]�Ͻ'�Ͻ�Ͻ��ϽߍϽ��Ͻ��Ͻ5�ϽX�Ͻ߁Ͻx�Ͻ�Ͻz�Ͻ<�Ͻ��ϽȊϽP   P   ��Ͻ��Ͻ��ϽR�Ͻ&�ϽE�ϽB�Ͻ��Ͻ��Ͻn�ϽI�ϽˈϽ5�ϽׂϽ�ϽϽقϽ5�Ͻ�Ͻx�ϽP   P   ��Ͻ��Ͻ��Ͻ�Ͻ}�Ͻ�Ͻ]�Ͻ��ϽʖϽ��ϽÏϽI�Ͻ��Ͻj�Ͻ؂Ͻ��Ͻ��Ͻz�Ͻ��ϽS�ϽP   P   ��ϽܓϽ�Ͻ��Ͻ@�Ͻ�Ͻ�Ͻo�Ͻ��Ͻ�Ͻ��Ͻn�Ͻ��ϽG�Ͻ��Ͻ�Ͻ�Ͻo�Ͻk�ϽʊϽP   P   �Ͻ��Ͻ��Ͻ��ϽC�Ͻg�Ͻ�ϽS�Ͻ�Ͻ��ϽʖϽ��ϽߍϽ�ϽϽF�Ͻ\�Ͻo�ϽφϽ�ϽP   P   ��Ͻ��ϽҕϽ�ϽN�ϽR�Ͻ��Ͻ��ϽS�Ͻo�Ͻ��Ͻ��Ͻ��Ͻ��ϽE�Ͻ��Ͻ��Ͻ`�Ͻ��Ͻ-�ϽP   P   �Ͻ��Ͻ�Ͻ4�Ͻ|�Ͻ�Ͻ(�Ͻ��Ͻ�Ͻ�Ͻ]�ϽB�Ͻ�Ͻ��ϽމϽ��ϽфϽ̃Ͻ�Ͻ��ϽP   P   ��Ͻ�Ͻ��ϽR�Ͻ0�Ͻ��Ͻ�ϽR�Ͻg�Ͻ�Ͻ�ϽE�Ͻ'�Ͻ��Ͻ6�Ͻ��ϽN�Ͻ��Ͻ݃Ͻ1�ϽP   P   ��ϽD�Ͻ6�ϽZ�Ͻj�Ͻ0�Ͻ|�ϽN�ϽC�Ͻ@�Ͻ}�Ͻ&�Ͻ]�Ͻw�Ͻ'�Ͻ,�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   �Ͻh�Ͻ�ϽʌϽZ�ϽR�Ͻ4�Ͻ�Ͻ��Ͻ��Ͻ�ϽR�ϽM�Ͻs�ϽȌϽ�Ͻ��Ͻ�ϽفϽ́ϽP   P   t�Ͻ�ϽF�Ͻ�Ͻ6�Ͻ��Ͻ�ϽҕϽ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ'�Ͻ�Ͻ�Ͻ�Ͻ~�Ͻ��ϽP   P   ��ϽP�Ͻ�Ͻh�ϽD�Ͻ�Ͻ��Ͻ��Ͻ��ϽܓϽ��Ͻ��Ͻ��Ͻ֍Ͻ4�ϽK�Ͻ��ϽK�Ͻo�Ͻ��ϽP   P   ʄϽ��Ͻ��Ͻ܇Ͻ�Ͻ �Ͻ�Ͻ��Ͻ;�Ͻ��Ͻ��ϽڏϽ\�Ͻ؎Ͻ(�Ͻ��Ͻw�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ[�Ͻ�Ͻ�ϽH�Ͻ��Ͻ!�Ͻ��Ͻ��Ͻ��ϽS�Ͻ΍ϽՌϽΌϽ��Ͻ*�ϽЈϽ
�Ͻ	�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ�Ͻ,�ϽчϽ��Ͻ��Ͻ�Ͻ��ϽϽ{�Ͻ��Ͻ؊Ͻ7�Ͻ��Ͻ҈ϽƇϽ��Ͻ	�ϽP   P   ��ϽR�ϽW�Ͻ��Ͻ]�Ͻ��Ͻ�Ͻj�ϽY�ϽΈϽ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻp�Ͻ��ϽƇϽ
�ϽP   P   w�Ͻ^�ϽȈϽ��Ͻ�Ͻ҈Ͻ��Ͻ��Ͻa�ϽG�Ͻ��Ͻ|�ϽׇϽ��Ͻ��ϽA�Ͻ��Ͻp�Ͻ҈ϽЈϽP   P   ��Ͻ(�ϽǋϽ��ϽZ�Ͻ�Ͻ;�Ͻu�Ͻ[�ϽE�Ͻ��Ͻ��Ͻ9�Ͻ(�Ͻ{�Ͻ�ϽA�Ͻ��Ͻ��Ͻ*�ϽP   P   )�Ͻ׍Ͻk�ϽՍϽ)�ϽԍϽ�Ͻ��Ͻ�Ͻ��Ͻo�Ͻ��Ͻh�Ͻ��Ͻ��Ͻ{�Ͻ��Ͻ��Ͻ7�Ͻ��ϽP   P   ؎Ͻ��Ͻ��ϽT�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ̊Ͻr�Ͻ��Ͻ-�Ͻ��Ͻ��Ͻ(�Ͻ��Ͻ��Ͻ؊ϽΌϽP   P   \�Ͻh�Ͻ)�ϽΓϽ��Ͻ��Ͻ�Ͻ��Ͻ%�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ-�Ͻh�Ͻ9�ϽׇϽ�Ͻ��ϽՌϽP   P   ڏϽ3�Ͻ��Ͻa�Ͻ8�ϽG�Ͻ��Ͻ͔Ͻ�ϽɏϽ��ϽP�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ|�Ͻ�Ͻ{�Ͻ΍ϽP   P   ��ϽӒϽΕϽ�Ͻ}�Ͻ��ϽT�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻr�Ͻo�Ͻ��Ͻ��Ͻ��ϽϽS�ϽP   P   ��Ͻ�Ͻ��ϽX�ϽҚϽt�Ͻ��Ͻ�ϽJ�Ͻ��Ͻ�ϽɏϽ�Ͻ̊Ͻ��ϽE�ϽG�ϽΈϽ��Ͻ��ϽP   P   ;�ϽБϽɕϽ-�Ͻy�Ͻ��Ͻ~�Ͻ��ϽV�ϽJ�Ͻ��Ͻ�Ͻ%�Ͻ��Ͻ�Ͻ[�Ͻa�ϽY�Ͻ�Ͻ��ϽP   P   ��Ͻ��Ͻ�Ͻ�Ͻ̚Ͻ؜Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ͔Ͻ��Ͻ��Ͻ��Ͻu�Ͻ��Ͻj�Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻ�ϽE�Ͻs�Ͻ��Ͻl�Ͻ��Ͻ~�Ͻ��ϽT�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ;�Ͻ��Ͻ�Ͻ��Ͻ!�ϽP   P    �Ͻ��Ͻ��Ͻ��Ͻ:�Ͻ��Ͻ��Ͻ؜Ͻ��Ͻt�Ͻ��ϽG�Ͻ��Ͻ��ϽԍϽ�Ͻ҈Ͻ��ϽчϽ��ϽP   P   �ϽQ�ϽK�Ͻi�ϽϽ:�Ͻs�Ͻ̚Ͻy�ϽҚϽ}�Ͻ8�Ͻ��Ͻ��Ͻ)�ϽZ�Ͻ�Ͻ]�Ͻ,�ϽH�ϽP   P   ܇ϽR�Ͻ��Ͻ�Ͻi�Ͻ��ϽE�Ͻ�Ͻ-�ϽX�Ͻ�Ͻa�ϽΓϽT�ϽՍϽ��Ͻ��Ͻ��Ͻ�Ͻ�ϽP   P   ��ϽU�ϽֈϽ��ϽK�Ͻ��Ͻ�Ͻ�ϽɕϽ��ϽΕϽ��Ͻ)�Ͻ��Ͻk�ϽǋϽȈϽW�Ͻ��Ͻ�ϽP   P   ��Ͻ��ϽU�ϽR�ϽQ�Ͻ��Ͻ��Ͻ��ϽБϽ�ϽӒϽ3�Ͻh�Ͻ��Ͻ׍Ͻ(�Ͻ^�ϽR�Ͻ��Ͻ[�ϽP   P   �Ͻ��ϽԉϽ7�Ͻ7�Ͻ��Ͻ\�Ͻ��Ͻ�Ͻ�Ͻ<�Ͻ��ϽA�Ͻ܏Ͻ��Ͻt�Ͻ��ϽJ�Ͻ��ϽʉϽP   P   ʉϽ��Ͻ��Ͻb�Ͻ=�Ͻw�Ͻ�Ͻ��ϽU�Ͻ؏Ͻ��Ͻ�Ͻ��Ͻ+�Ͻl�Ͻ�Ͻs�Ͻ�Ͻf�Ͻ��ϽP   P   ��Ͻ�Ͻ݉Ͻl�Ͻ�ϽċϽɋϽ��Ͻ��Ͻ��Ͻ$�ϽԍϽ$�Ͻ�ϽӌϽ�Ͻ�ϽˋϽ^�Ͻf�ϽP   P   J�Ͻ/�Ͻ]�Ͻ5�Ͻ8�ϽËϽ��Ͻ��Ͻ�Ͻo�Ͻ,�Ͻ��ϽˋϽ8�Ͻ4�Ͻ��Ͻ��Ͻ��ϽˋϽ�ϽP   P   ��Ͻx�Ͻ��Ͻ��ϽI�Ͻa�ϽǋϽ��Ͻ��Ͻy�ϽǊϽ��Ͻ(�ϽЊϽ	�Ͻb�Ͻ �Ͻ��Ͻ�Ͻs�ϽP   P   t�Ͻw�ϽL�Ͻ	�ϽҍϽz�Ͻ��Ͻu�Ͻ��Ͻ��Ͻ��Ͻ��ϽN�Ͻ:�Ͻa�ϽˊϽb�Ͻ��Ͻ�Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻ}�Ͻ\�Ͻl�Ͻb�Ͻ}�Ͻ��Ͻ5�Ͻ�Ͻp�Ͻ
�Ͻ�Ͻ��Ͻa�Ͻ	�Ͻ4�ϽӌϽl�ϽP   P   ܏Ͻ�Ͻ2�Ͻu�Ͻ͒Ͻ!�Ͻ�Ͻ��Ͻ/�Ͻ�Ͻ�Ͻ֊Ͻ?�Ͻ��Ͻ�Ͻ:�ϽЊϽ8�Ͻ�Ͻ+�ϽP   P   A�Ͻ?�Ͻ��ϽՔϽ�Ͻ��Ͻt�ϽZ�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ?�Ͻ
�ϽN�Ͻ(�ϽˋϽ$�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ֕ϽۖϽҖϽ
�Ͻ{�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ֊Ͻp�Ͻ��Ͻ��Ͻ��ϽԍϽ�ϽP   P   <�Ͻ�Ͻ:�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ	�Ͻ>�Ͻ!�Ͻ�Ͻ�Ͻ�Ͻ�Ͻ�Ͻ��ϽǊϽ,�Ͻ$�Ͻ��ϽP   P   �Ͻ �Ͻh�ϽɗϽ��Ͻ(�ϽM�Ͻ��ϽΗϽF�Ͻ!�Ͻ��Ͻ��Ͻ�Ͻ5�Ͻ��Ͻy�Ͻo�Ͻ��Ͻ؏ϽP   P   �ϽדϽH�ϽƗϽt�Ͻ��Ͻ��Ͻ՚Ͻg�ϽΗϽ>�Ͻ�Ͻ�Ͻ/�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽU�ϽP   P   ��Ͻ��ϽǔϽ�Ͻ��Ͻ͚Ͻ͛Ͻ��Ͻ՚Ͻ��Ͻ	�Ͻ{�ϽZ�Ͻ��Ͻ}�Ͻu�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   \�Ͻ�Ͻ*�ϽەϽ��ϽM�ϽV�Ͻ͛Ͻ��ϽM�Ͻ��Ͻ
�Ͻt�Ͻ�Ͻb�Ͻ��ϽǋϽ��ϽɋϽ�ϽP   P   ��Ͻq�Ͻ(�Ͻ��Ͻ��Ͻ{�ϽM�Ͻ͚Ͻ��Ͻ(�Ͻ��ϽҖϽ��Ͻ!�Ͻl�Ͻz�Ͻa�ϽËϽċϽw�ϽP   P   7�Ͻ��Ͻ?�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻt�Ͻ��Ͻ��ϽۖϽ�Ͻ͒Ͻ\�ϽҍϽI�Ͻ8�Ͻ�Ͻ=�ϽP   P   7�Ͻ��Ͻ-�Ͻ��Ͻ��Ͻ��ϽەϽ�ϽƗϽɗϽ�Ͻ֕ϽՔϽu�Ͻ}�Ͻ	�Ͻ��Ͻ5�Ͻl�Ͻb�ϽP   P   ԉϽL�Ͻz�Ͻ-�Ͻ?�Ͻ(�Ͻ*�ϽǔϽH�Ͻh�Ͻ:�Ͻ��Ͻ��Ͻ2�Ͻ��ϽL�Ͻ��Ͻ]�Ͻ݉Ͻ��ϽP   P   ��Ͻ�ϽL�Ͻ��Ͻ��Ͻq�Ͻ�Ͻ��ϽדϽ �Ͻ�Ͻ��Ͻ?�Ͻ�Ͻ��Ͻw�Ͻx�Ͻ/�Ͻ�Ͻ��ϽP   P   ��Ͻe�ϽڍϽ>�Ͻ�Ͻv�ϽI�Ͻ��Ͻ<�Ͻ�Ͻ��Ͻ��Ͻ}�Ͻ+�Ͻe�Ͻa�Ͻl�ϽM�Ͻ�Ͻd�ϽP   P   d�Ͻ��Ͻ�Ͻ;�Ͻ��Ͻ>�Ͻ%�Ͻ_�Ͻ��ϽF�ϽF�Ͻ#�ϽX�Ͻ��ϽP�Ͻ:�Ͻ$�Ͻ��Ͻ�Ͻ�ϽP   P   �Ͻ��ϽӍϽ	�Ͻ��Ͻ.�Ͻ֎Ͻr�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ$�Ͻ�Ͻ[�Ͻ��Ͻ��Ͻ@�Ͻ3�Ͻ�ϽP   P   M�Ͻ\�Ͻq�Ͻl�Ͻ��Ͻh�Ͻ�Ͻ�Ͻ]�Ͻ
�Ͻ��Ͻ`�Ͻk�Ͻ��Ͻ��ϽV�ϽގϽ�Ͻ@�Ͻ��ϽP   P   l�Ͻ#�Ͻ��Ͻ��Ͻ?�Ͻ�Ͻ�Ͻ��Ͻr�Ͻ��Ͻ�Ͻk�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽގϽ��Ͻ$�ϽP   P   a�Ͻ��Ͻ��Ͻ��Ͻ̐Ͻ��Ͻ!�Ͻ��Ͻo�Ͻ��Ͻ��Ͻ?�Ͻ׍Ͻ��Ͻ�Ͻ��Ͻ��ϽV�Ͻ��Ͻ:�ϽP   P   e�ϽڑϽ��Ͻ��Ͻ��Ͻ��Ͻp�Ͻ?�Ͻ0�ϽʎϽ��Ͻ�Ͻj�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ[�ϽP�ϽP   P   +�Ͻ�ϽђϽ��Ͻ��ϽےϽ'�Ͻ�Ͻ��Ͻ-�Ͻ��Ͻ��Ͻ��Ͻ2�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽP   P   }�ϽѓϽ�Ͻ�ϽI�Ͻ��Ͻ�Ͻ��Ͻx�Ͻ/�Ͻ�ϽV�Ͻv�Ͻ��Ͻj�Ͻ׍Ͻ��Ͻk�Ͻ$�ϽX�ϽP   P   ��Ͻ1�Ͻ�Ͻ��Ͻ_�Ͻn�Ͻ��ϽĕϽF�Ͻ��Ͻ/�ϽÐϽV�Ͻ��Ͻ�Ͻ?�Ͻk�Ͻ`�Ͻ��Ͻ#�ϽP   P   ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻx�Ͻ	�Ͻ��Ͻ&�ϽДϽ��Ͻ/�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�ϽF�ϽP   P   �ϽĔϽ��ϽɗϽ��Ͻ1�ϽX�ϽݘϽ�Ͻ��ϽДϽ��Ͻ/�Ͻ-�ϽʎϽ��Ͻ��Ͻ
�Ͻ��ϽF�ϽP   P   <�ϽU�Ͻ
�Ͻ��Ͻ��Ͻ'�Ͻ$�Ͻ!�Ͻ��Ͻ�Ͻ&�ϽF�Ͻx�Ͻ��Ͻ0�Ͻo�Ͻr�Ͻ]�Ͻ�Ͻ��ϽP   P   ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ �Ͻ��ϽP�Ͻ!�ϽݘϽ��ϽĕϽ��Ͻ�Ͻ?�Ͻ��Ͻ��Ͻ�Ͻr�Ͻ_�ϽP   P   I�ϽP�Ͻ��Ͻ��Ͻ��Ͻ{�Ͻ�Ͻ��Ͻ$�ϽX�Ͻ	�Ͻ��Ͻ�Ͻ&�Ͻp�Ͻ!�Ͻ�Ͻ�Ͻ֎Ͻ%�ϽP   P   v�ϽʑϽ�Ͻ�Ͻ��Ͻ;�Ͻ{�Ͻ �Ͻ'�Ͻ1�Ͻx�Ͻn�Ͻ��ϽےϽ��Ͻ��Ͻ�Ͻh�Ͻ.�Ͻ>�ϽP   P   �Ͻ��Ͻ��Ͻ̓Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ_�ϽI�Ͻ��Ͻ��Ͻ̐Ͻ?�Ͻ��Ͻ��Ͻ��ϽP   P   >�ϽR�Ͻ��Ͻ�Ͻ̓Ͻ�Ͻ��Ͻ��Ͻ��ϽɗϽ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻl�Ͻ	�Ͻ;�ϽP   P   ڍϽi�ϽQ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ
�Ͻ��Ͻ�Ͻ�Ͻ�ϽђϽ��Ͻ��Ͻ��Ͻq�ϽӍϽ�ϽP   P   e�Ͻ��Ͻi�ϽR�Ͻ��ϽʑϽP�Ͻ�ϽU�ϽĔϽ�Ͻ1�ϽѓϽ�ϽڑϽ��Ͻ#�Ͻ\�Ͻ��Ͻ��ϽP   P   O�ϽR�ϽӐϽk�ϽƑϽV�Ͻ�Ͻ��Ͻ��Ͻ�Ͻb�Ͻ�Ͻ��Ͻ��Ͻ�ϽS�ϽđϽ_�Ͻ�Ͻ[�ϽP   P   [�Ͻ��ϽE�ϽِϽ��ϽÑϽ-�Ͻ�Ͻ
�Ͻ��Ͻ�ϽÓϽ��Ͻ��Ͻ3�Ͻ9�Ͻ��Ͻ�Ͻ��ϽK�ϽP   P   �Ͻ��Ͻ�Ͻ��Ͻ>�Ͻo�ϽȑϽ��Ͻ�Ͻ̒Ͻ��Ͻ��Ͻ�Ͻ�Ͻ �Ͻ��Ͻ̑Ͻ��Ͻ6�Ͻ��ϽP   P   _�ϽL�Ͻ^�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽC�Ͻ��Ͻ�Ͻ
�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   đϽ
�Ͻ��ϽבϽ�Ͻ��ϽΑϽޑϽÑϽs�Ͻ��ϽL�Ͻ��ϽV�Ͻ��Ͻ��ϽɑϽ��Ͻ̑Ͻ��ϽP   P   S�ϽG�Ͻ�Ͻ�Ͻ7�Ͻa�Ͻ�Ͻ��Ͻ��Ͻz�Ͻ��Ͻ��ϽِϽĐϽȐϽ̐Ͻ��Ͻ��Ͻ��Ͻ9�ϽP   P   �Ͻ��Ͻ#�Ͻ	�Ͻ6�Ͻ��Ͻ-�Ͻ�Ͻ!�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽȐϽ��Ͻ�Ͻ �Ͻ3�ϽP   P   ��Ͻ��Ͻ�Ͻp�Ͻ-�Ͻ.�Ͻ��Ͻ��Ͻ�ϽؒϽ%�ϽV�ϽѐϽ�Ͻ�ϽĐϽV�Ͻ
�Ͻ�Ͻ��ϽP   P   ��Ͻn�Ͻ͕Ͻ|�Ͻ��Ͻy�Ͻ��Ͻ<�Ͻ�Ͻ��ϽҒϽ��Ͻ�ϽѐϽ��ϽِϽ��Ͻ�Ͻ�Ͻ��ϽP   P   �Ͻs�Ͻx�ϽJ�Ͻ	�Ͻ�Ͻ(�Ͻ��Ͻ��ϽݔϽ͓Ͻ��Ͻ��ϽV�Ͻ��Ͻ��ϽL�Ͻ��Ͻ��ϽÓϽP   P   b�Ͻ	�ϽB�Ͻ��Ͻ[�ϽJ�ϽX�Ͻ�Ͻ'�Ͻ�Ͻ��Ͻ͓ϽҒϽ%�Ͻ��Ͻ��Ͻ��ϽC�Ͻ��Ͻ�ϽP   P   �Ͻ�Ͻ��Ͻ��Ͻ��Ͻk�Ͻx�Ͻ��Ͻ��Ͻ�Ͻ�ϽݔϽ��ϽؒϽ�Ͻz�Ͻs�Ͻ�Ͻ̒Ͻ��ϽP   P   ��ϽĕϽ.�ϽژϽ�Ͻ�Ͻ�Ͻ�Ͻ�Ͻ��Ͻ'�Ͻ��Ͻ�Ͻ�Ͻ!�Ͻ��ϽÑϽ��Ͻ�Ͻ
�ϽP   P   ��ϽK�Ͻo�Ͻ�Ͻ��Ͻ��Ͻh�ϽO�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ<�Ͻ��Ͻ�Ͻ��ϽޑϽ��Ͻ��Ͻ�ϽP   P   �Ͻ��Ͻ��Ͻq�Ͻ9�Ͻ��Ͻ�Ͻh�Ͻ�Ͻx�ϽX�Ͻ(�Ͻ��Ͻ��Ͻ-�Ͻ�ϽΑϽ��ϽȑϽ-�ϽP   P   V�ϽۓϽ�ϽT�Ͻ�Ͻ?�Ͻ��Ͻ��Ͻ�Ͻk�ϽJ�Ͻ�Ͻy�Ͻ.�Ͻ��Ͻa�Ͻ��Ͻ��Ͻo�ϽÑϽP   P   ƑϽ(�Ͻ*�Ͻa�Ͻ~�Ͻ�Ͻ9�Ͻ��Ͻ�Ͻ��Ͻ[�Ͻ	�Ͻ��Ͻ-�Ͻ6�Ͻ7�Ͻ�Ͻ��Ͻ>�Ͻ��ϽP   P   k�Ͻ�Ͻ�Ͻ�Ͻa�ϽT�Ͻq�Ͻ�ϽژϽ��Ͻ��ϽJ�Ͻ|�Ͻp�Ͻ	�Ͻ�ϽבϽ��Ͻ��ϽِϽP   P   ӐϽE�ϽёϽ�Ͻ*�Ͻ�Ͻ��Ͻo�Ͻ.�Ͻ��ϽB�Ͻx�Ͻ͕Ͻ�Ͻ#�Ͻ�Ͻ��Ͻ^�Ͻ�ϽE�ϽP   P   R�Ͻ��ϽE�Ͻ�Ͻ(�ϽۓϽ��ϽK�ϽĕϽ�Ͻ	�Ͻs�Ͻn�Ͻ��Ͻ��ϽG�Ͻ
�ϽL�Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻ�Ͻ��Ͻ.�Ͻ�Ͻo�ϽҖϽP�Ͻ��Ͻ��Ͻ��ϽV�Ͻ��Ͻ=�Ͻg�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��ϽٓϽ��Ͻ��Ͻ9�Ͻa�Ͻ2�Ͻ��Ͻ�ϽݕϽ��Ͻm�Ͻ��ϽO�Ͻ��Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ|�Ͻ��Ͻ��Ͻ��Ͻp�Ͻn�Ͻ�Ͻ�Ͻ̔Ͻ(�ϽϔϽ,�Ͻ��Ͻ�Ͻ�ϽU�ϽY�ϽÓϽ�ϽP   P   ��Ͻ	�Ͻ�Ͻ��ϽʓϽL�Ͻ��Ͻ��ϽҔϽ�Ͻ�Ͻx�Ͻ��Ͻ�Ͻ$�Ͻ��ϽݓϽʓϽY�Ͻ��ϽP   P   g�ϽݔϽ��Ͻ��Ͻ��ϽÔϽb�Ͻ�Ͻ�Ͻ��ϽÓϽ��Ͻ5�ϽœϽƓϽ�Ͻ�ϽݓϽU�Ͻ��ϽP   P   =�Ͻ�Ͻ
�Ͻ<�ϽݔϽ)�ϽE�ϽՔϽ˔Ͻ�ϽB�ϽГϽ��ϽݓϽ�Ͻ�Ͻ�Ͻ��Ͻ�ϽO�ϽP   P   ��Ͻh�ϽԕϽF�Ͻ֕Ͻc�Ͻ�Ͻ��Ͻ�ϽI�Ͻ��Ͻ��Ͻ��ϽS�Ͻ~�Ͻ�ϽƓϽ$�Ͻ�Ͻ��ϽP   P   V�Ͻ0�Ͻ	�Ͻ�ϽʖϽ/�Ͻ3�ϽD�ϽR�Ͻ��Ͻ.�ϽʓϽÓϽ�ϽS�ϽݓϽœϽ�Ͻ��Ͻm�ϽP   P   ��Ͻ�Ͻ-�Ͻ��Ͻi�Ͻ��Ͻ��ϽܖϽ��Ͻ��Ͻ$�Ͻy�Ͻ9�ϽÓϽ��Ͻ��Ͻ5�Ͻ��Ͻ,�Ͻ��ϽP   P   ��ϽЗϽ�Ͻo�Ͻs�Ͻw�ϽB�Ͻ^�ϽŗϽo�Ͻ�ϽܔϽy�ϽʓϽ��ϽГϽ��Ͻx�ϽϔϽݕϽP   P   ��Ͻ=�ϽV�ϽۘϽI�Ͻ��ϽO�Ͻ�Ͻ�Ͻ_�Ͻ�Ͻ�Ͻ$�Ͻ.�Ͻ��ϽB�ϽÓϽ�Ͻ(�Ͻ�ϽP   P   P�Ͻw�Ͻy�Ͻ��ϽP�ϽC�Ͻ+�ϽR�Ͻ��Ͻ��Ͻ_�Ͻo�Ͻ��Ͻ��ϽI�Ͻ�Ͻ��Ͻ�Ͻ̔Ͻ��ϽP   P   ҖϽڗϽ5�Ͻc�Ͻ��Ͻ��Ͻc�Ͻv�Ͻ��Ͻ��Ͻ�ϽŗϽ��ϽR�Ͻ�Ͻ˔Ͻ�ϽҔϽ�Ͻ2�ϽP   P   o�ϽŖϽ�Ͻ�ϽW�Ͻ��Ͻ��Ͻ��Ͻv�ϽR�Ͻ�Ͻ^�ϽܖϽD�Ͻ��ϽՔϽ�Ͻ��Ͻ�Ͻa�ϽP   P   �Ͻ�Ͻ{�Ͻe�Ͻ.�Ͻ�Ͻ��Ͻ��Ͻc�Ͻ+�ϽO�ϽB�Ͻ��Ͻ3�Ͻ�ϽE�Ͻb�Ͻ��Ͻn�Ͻ9�ϽP   P   .�Ͻ]�Ͻ�Ͻ��Ͻ]�Ͻ�Ͻ�Ͻ��Ͻ��ϽC�Ͻ��Ͻw�Ͻ��Ͻ/�Ͻc�Ͻ)�ϽÔϽL�Ͻp�Ͻ��ϽP   P   ��Ͻ��Ͻ�Ͻ�Ͻ˗Ͻ]�Ͻ.�ϽW�Ͻ��ϽP�ϽI�Ͻs�Ͻi�ϽʖϽ֕ϽݔϽ��ϽʓϽ��Ͻ��ϽP   P   �Ͻ��Ͻ �Ͻ��Ͻ�Ͻ��Ͻe�Ͻ�Ͻc�Ͻ��ϽۘϽo�Ͻ��Ͻ�ϽF�Ͻ<�Ͻ��Ͻ��Ͻ��ϽٓϽP   P   ��Ͻ�Ͻ��Ͻ �Ͻ�Ͻ�Ͻ{�Ͻ�Ͻ5�Ͻy�ϽV�Ͻ�Ͻ-�Ͻ	�ϽԕϽ
�Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ]�Ͻ�ϽŖϽڗϽw�Ͻ=�ϽЗϽ�Ͻ0�Ͻh�Ͻ�ϽݔϽ	�Ͻ|�Ͻ��ϽP   P   O�Ͻ�ϽN�Ͻ��ϽW�Ͻ^�Ͻ��Ͻ�ϽחϽ>�Ͻ�Ͻ��Ͻ��Ͻ�Ͻl�Ͻs�Ͻ��Ͻx�Ͻ?�Ͻ�ϽP   P   �Ͻ��ϽY�Ͻ~�ϽB�Ͻa�Ͻe�Ͻ@�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ&�ϽG�Ͻ}�Ͻ��Ͻy�Ͻ��Ͻ(�ϽP   P   ?�Ͻ��ϽN�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ7�Ͻ��ϽG�Ͻ�ϽU�Ͻu�Ͻ�Ͻ~�Ͻ��Ͻ��ϽQ�Ͻ��ϽP   P   x�Ͻk�Ͻ��Ͻf�Ͻu�ϽV�Ͻ2�Ͻ��Ͻw�ϽіϽ��Ͻ#�Ͻ�Ͻ7�ϽؖϽ��Ͻ	�Ͻ]�Ͻ��Ͻy�ϽP   P   ��Ͻ�Ͻ˖Ͻ�Ͻ�Ͻ��ϽϖϽ1�Ͻ��Ͻ��Ͻ�Ͻ��Ͻk�Ͻ��Ͻ�Ͻ��Ͻa�Ͻ	�Ͻ��Ͻ��ϽP   P   s�Ͻ��Ͻp�Ͻ�Ͻ��ϽU�Ͻ��ϽP�Ͻc�Ͻv�Ͻ��Ͻ �Ͻ�ϽS�Ͻ=�Ͻ��Ͻ��Ͻ��Ͻ~�Ͻ}�ϽP   P   l�Ͻ��Ͻ�ϽE�ϽԗϽ�ϽZ�Ͻ[�Ͻ�Ͻ�Ͻ͖ϽK�ϽO�Ͻ*�Ͻ�Ͻ=�Ͻ�ϽؖϽ�ϽG�ϽP   P   �Ͻ��Ͻ��Ͻ��ϽV�Ͻ��Ͻ|�Ͻ��Ͻ�Ͻ0�Ͻ,�Ͻ��Ͻ8�Ͻ�Ͻ*�ϽS�Ͻ��Ͻ7�Ͻu�Ͻ&�ϽP   P   ��Ͻc�ϽN�Ͻ�Ͻ��Ͻ?�Ͻ�Ͻ��Ͻs�ϽЗϽD�Ͻ�Ͻ�Ͻ8�ϽO�Ͻ�Ͻk�Ͻ�ϽU�Ͻ��ϽP   P   ��ϽԘϽ��Ͻ�ϽV�ϽG�Ͻ��Ͻ͙Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��ϽK�Ͻ �Ͻ��Ͻ#�Ͻ�Ͻ�ϽP   P   �ϽB�Ͻz�Ͻ	�Ͻy�Ͻ��Ͻ��Ͻ3�Ͻ8�Ͻ��Ͻ��Ͻ�ϽD�Ͻ,�Ͻ͖Ͻ��Ͻ�Ͻ��ϽG�Ͻ��ϽP   P   >�Ͻ��Ͻ�ϽܚϽΚϽ�Ͻ̚ϽۚϽ��Ͻ�Ͻ��Ͻ��ϽЗϽ0�Ͻ�Ͻv�Ͻ��ϽіϽ��Ͻ��ϽP   P   חϽ��Ͻ��Ͻ��Ͻ2�Ͻ��Ͻ-�Ͻ��Ͻ:�Ͻ��Ͻ8�Ͻ��Ͻs�Ͻ�Ͻ�Ͻc�Ͻ��Ͻw�Ͻ7�Ͻ��ϽP   P   �ϽM�Ͻ|�Ͻa�Ͻ֚Ͻ�Ͻ��ϽϽ��ϽۚϽ3�Ͻ͙Ͻ��Ͻ��Ͻ[�ϽP�Ͻ1�Ͻ��Ͻ��Ͻ@�ϽP   P   ��Ͻ9�Ͻ��ϽșϽ��Ͻ��Ͻ>�Ͻ��Ͻ-�Ͻ̚Ͻ��Ͻ��Ͻ�Ͻ|�ϽZ�Ͻ��ϽϖϽ2�Ͻ��Ͻe�ϽP   P   ^�Ͻ��Ͻ��Ͻ�Ͻ"�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��ϽG�Ͻ?�Ͻ��Ͻ�ϽU�Ͻ��ϽV�Ͻ��Ͻa�ϽP   P   W�Ͻ��Ͻ-�ϽS�Ͻ��Ͻ"�Ͻ��Ͻ֚Ͻ2�ϽΚϽy�ϽV�Ͻ��ϽV�ϽԗϽ��Ͻ�Ͻu�Ͻ��ϽB�ϽP   P   ��Ͻ��Ͻ��Ͻ�ϽS�Ͻ�ϽșϽa�Ͻ��ϽܚϽ	�Ͻ�Ͻ�Ͻ��ϽE�Ͻ�Ͻ�Ͻf�Ͻ��Ͻ~�ϽP   P   N�Ͻ{�Ͻ%�Ͻ��Ͻ-�Ͻ��Ͻ��Ͻ|�Ͻ��Ͻ�Ͻz�Ͻ��ϽN�Ͻ��Ͻ�Ͻp�Ͻ˖Ͻ��ϽN�ϽY�ϽP   P   �ϽM�Ͻ{�Ͻ��Ͻ��Ͻ��Ͻ9�ϽM�Ͻ��Ͻ��ϽB�ϽԘϽc�Ͻ��Ͻ��Ͻ��Ͻ�Ͻk�Ͻ��Ͻ��ϽP   P   �Ͻ�Ͻ��Ͻ�Ͻ(�Ͻa�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ,�Ͻ��Ͻ��Ͻ�Ͻ�Ͻm�Ͻ�Ͻ�Ͻ��Ͻ�ϽP   P   �Ͻ�Ͻj�Ͻt�Ͻi�ϽI�ϽҙϽ��Ͻ��Ͻ�Ͻ�ϽԙϽ��Ͻ��Ͻ��Ͻ��Ͻb�Ͻ{�Ͻ��Ͻa�ϽP   P   ��Ͻ�Ͻ��Ͻ_�Ͻ�Ͻ�Ͻs�Ͻ��Ͻ0�Ͻ_�ϽR�Ͻ��ϽN�ϽG�Ͻ�ϽÙϽ:�Ͻ��Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻo�Ͻ��Ͻ	�Ͻ�ϽژϽ�Ͻ��Ͻ�Ͻ/�Ͻ%�Ͻ�Ͻ��Ͻ��Ͻ{�ϽP   P   �Ͻ�ϽT�Ͻ(�Ͻ�ϽE�Ͻf�Ͻ�ϽX�Ͻ+�Ͻ�Ͻ�Ͻ~�ϽјϽ�Ͻ*�Ͻ3�Ͻ�Ͻ:�Ͻb�ϽP   P   m�Ͻ��Ͻ��Ͻ��Ͻf�Ͻc�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ]�Ͻ��ϽߘϽ�Ͻ��Ͻd�Ͻ*�Ͻ%�ϽÙϽ��ϽP   P   �Ͻ�Ͻ��Ͻ'�Ͻ�Ͻ#�Ͻ|�Ͻ~�Ͻ?�Ͻ<�Ͻ��Ͻ��ϽޘϽ�Ͻ��Ͻ��Ͻ�Ͻ/�Ͻ�Ͻ��ϽP   P   �Ͻi�Ͻ:�ϽǚϽ��Ͻ/�Ͻ?�Ͻ��Ͻ��Ͻ)�Ͻ�Ͻ��Ͻ�ϽޘϽ�Ͻ�ϽјϽ�ϽG�Ͻ��ϽP   P   ��ϽޚϽ��ϽКϽW�Ͻ�Ͻ��Ͻ��Ͻs�Ͻ�Ͻm�Ͻ��Ͻ��Ͻ�ϽޘϽߘϽ~�Ͻ��ϽN�Ͻ��ϽP   P   ��Ͻ
�Ͻ��Ͻ4�Ͻ+�Ͻ �Ͻ�Ͻ�Ͻ�Ͻ��ϽҙϽ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��ϽԙϽP   P   ,�Ͻ��Ͻ1�Ͻ��Ͻ��Ͻ4�ϽÛϽ��ϽN�Ͻ��Ͻ��ϽҙϽm�Ͻ�Ͻ��Ͻ]�Ͻ�ϽژϽR�Ͻ�ϽP   P   ��Ͻ��Ͻ�Ͻ��Ͻe�Ͻt�Ͻ[�ϽN�ϽڛϽ�Ͻ��Ͻ��Ͻ�Ͻ)�Ͻ<�Ͻ�Ͻ+�Ͻ�Ͻ_�Ͻ�ϽP   P   ��Ͻ��ϽB�ϽӛϽ�Ͻ��Ͻ�Ͻ��Ͻ�ϽڛϽN�Ͻ�Ͻs�Ͻ��Ͻ?�Ͻ�ϽX�Ͻ	�Ͻ0�Ͻ��ϽP   P   ��ϽܚϽۚϽ��ϽO�Ͻ˜Ͻq�Ͻ��Ͻ��ϽN�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ~�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ<�ϽךϽ �Ͻ��ϽS�Ͻ�Ͻq�Ͻ�Ͻ[�ϽÛϽ�Ͻ��Ͻ?�Ͻ|�Ͻ��Ͻf�Ͻo�Ͻs�ϽҙϽP   P   a�Ͻ��Ͻ6�ϽȚϽ�ϽI�ϽS�Ͻ˜Ͻ��Ͻt�Ͻ4�Ͻ �Ͻ�Ͻ/�Ͻ#�Ͻc�ϽE�Ͻ�Ͻ�ϽI�ϽP   P   (�Ͻm�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��ϽO�Ͻ�Ͻe�Ͻ��Ͻ+�ϽW�Ͻ��Ͻ�Ͻf�Ͻ�Ͻ��Ͻ�Ͻi�ϽP   P   �Ͻ��Ͻ��Ͻ�Ͻ��ϽȚϽ �Ͻ��ϽӛϽ��Ͻ��Ͻ4�ϽКϽǚϽ'�Ͻ��Ͻ(�Ͻ�Ͻ_�Ͻt�ϽP   P   ��Ͻ��Ͻq�Ͻ��Ͻ�Ͻ6�ϽךϽۚϽB�Ͻ�Ͻ1�Ͻ��Ͻ��Ͻ:�Ͻ��Ͻ��ϽT�Ͻ�Ͻ��Ͻj�ϽP   P   �ϽؘϽ��Ͻ��Ͻm�Ͻ��Ͻ<�ϽܚϽ��Ͻ��Ͻ��Ͻ
�ϽޚϽi�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�ϽP   P   ��Ͻ��Ͻ4�ϽB�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�Ͻ7�Ͻ�Ͻ�Ͻ'�Ͻ��Ͻ��ϽO�ϽW�Ͻ=�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻl�Ͻ�ϽQ�Ͻ��Ͻ֛Ͻ��ϽɛϽ��Ͻ�Ͻ�Ͻ}�ϽƛϽ��Ͻ7�Ͻ�ϽC�Ͻ��ϽP   P   =�Ͻ��Ͻm�Ͻ.�Ͻ�ϽP�Ͻ�Ͻ_�Ͻ��Ͻ͛ϽěϽ�Ͻ̛Ͻ͛ϽΛϽ_�Ͻ�Ͻs�Ͻ��ϽC�ϽP   P   W�ϽJ�Ͻ�ϽT�Ͻ�Ͻ��Ͻu�Ͻ+�Ͻc�Ͻ}�Ͻt�Ͻ��Ͻ��Ͻ`�Ͻ��Ͻ?�Ͻ�Ͻ}�Ͻs�Ͻ�ϽP   P   O�Ͻ��Ͻ��Ͻ��Ͻj�Ͻ	�Ͻ�Ͻ��Ͻ+�Ͻ0�Ͻ!�Ͻx�Ͻ��Ͻ��Ͻ�Ͻ3�ϽD�Ͻ�Ͻ�Ͻ7�ϽP   P   ��ϽۛϽ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ`�Ͻl�Ͻ!�Ͻx�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ3�Ͻ?�Ͻ_�Ͻ��ϽP   P   ��Ͻ��Ͻ
�Ͻ��Ͻ�Ͻ��Ͻ#�Ͻ��Ͻ͛ϽM�ϽC�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽΛϽƛϽP   P   '�Ͻ�Ͻ\�Ͻ+�Ͻ(�ϽC�Ͻ�Ͻ&�Ͻ��ϽܛϽR�Ͻm�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ`�Ͻ͛Ͻ}�ϽP   P   �Ͻ;�Ͻ��Ͻ6�Ͻm�Ͻ�ϽɜϽF�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ̛Ͻ�ϽP   P   �Ͻi�Ͻ��ϽX�Ͻ�Ͻ�Ͻb�ϽR�ϽW�Ͻ�Ͻ�Ͻ��Ͻ��Ͻm�Ͻ��Ͻ��Ͻx�Ͻ��Ͻ�Ͻ�ϽP   P   7�Ͻ�Ͻ9�Ͻ��Ͻ��Ͻ�ϽНϽ��Ͻ��Ͻ��ϽO�Ͻ�Ͻ��ϽR�ϽC�Ͻx�Ͻ!�Ͻt�ϽěϽ��ϽP   P   �Ͻ��Ͻ�Ͻ�Ͻ��ϽM�Ͻe�ϽȝϽ�Ͻ��Ͻ��Ͻ�Ͻ��ϽܛϽM�Ͻ!�Ͻ0�Ͻ}�Ͻ͛ϽɛϽP   P   �Ͻ��ϽF�ϽJ�Ͻ��Ͻ�Ͻ]�Ͻ�ϽɝϽ�Ͻ��ϽW�Ͻ�Ͻ��Ͻ͛Ͻl�Ͻ+�Ͻc�Ͻ��Ͻ��ϽP   P   �ϽI�Ͻ��Ͻ��ϽҝϽ	�Ͻ|�ϽW�Ͻ�ϽȝϽ��ϽR�ϽF�Ͻ&�Ͻ��Ͻ`�Ͻ��Ͻ+�Ͻ_�Ͻ֛ϽP   P   ��Ͻ2�Ͻd�Ͻr�Ͻ��Ͻ��Ͻ5�Ͻ|�Ͻ]�Ͻe�ϽНϽb�ϽɜϽ�Ͻ#�Ͻ��Ͻ�Ͻu�Ͻ�Ͻ��ϽP   P   ��Ͻ��Ͻb�Ͻ4�Ͻ��Ͻ�Ͻ��Ͻ	�Ͻ�ϽM�Ͻ�Ͻ�Ͻ�ϽC�Ͻ��Ͻ��Ͻ	�Ͻ��ϽP�ϽQ�ϽP   P   �ϽϛϽ�Ͻ7�Ͻ*�Ͻ��Ͻ��ϽҝϽ��Ͻ��Ͻ��Ͻ�Ͻm�Ͻ(�Ͻ�Ͻ��Ͻj�Ͻ�Ͻ�Ͻ�ϽP   P   B�Ͻ͛ϽÛϽڛϽ7�Ͻ4�Ͻr�Ͻ��ϽJ�Ͻ�Ͻ��ϽX�Ͻ6�Ͻ+�Ͻ��Ͻ��Ͻ��ϽT�Ͻ.�Ͻl�ϽP   P   4�Ͻ0�Ͻ`�ϽÛϽ�Ͻb�Ͻd�Ͻ��ϽF�Ͻ�Ͻ9�Ͻ��Ͻ��Ͻ\�Ͻ
�Ͻ��Ͻ��Ͻ�Ͻm�Ͻ��ϽP   P   ��ϽǚϽ0�Ͻ͛ϽϛϽ��Ͻ2�ϽI�Ͻ��Ͻ��Ͻ�Ͻi�Ͻ;�Ͻ�Ͻ��ϽۛϽ��ϽJ�Ͻ��Ͻ��ϽP   P   &�Ͻa�Ͻ<�Ͻ)�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�Ͻv�Ͻ��Ͻ!�ϽS�Ͻ-�Ͻ�ϽӝϽ�Ͻ5�ϽJ�Ͻc�ϽP   P   c�ϽY�Ͻ�Ͻ��Ͻ��Ͻ�ϽS�Ͻ��Ͻ,�Ͻ�Ͻ�Ͻ)�Ͻ?�ϽӝϽ��ϽR�ϽҝϽ\�Ͻm�Ͻ�ϽP   P   J�Ͻ�Ͻp�Ͻh�Ͻ[�Ͻk�Ͻs�Ͻ�Ͻ|�Ͻ��Ͻ��ϽK�Ͻ��Ͻ��ϽٝϽz�ϽŝϽ��Ͻ��Ͻm�ϽP   P   5�Ͻ��Ͻ^�Ͻ&�Ͻk�Ͻ��ϽG�Ͻ-�Ͻ��Ͻ��ϽɝϽP�ϽN�ϽÝϽ��Ͻ[�Ͻ�Ͻ�Ͻ��Ͻ\�ϽP   P   �Ͻ~�Ͻg�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ؝Ͻz�Ͻ��Ͻ:�Ͻ�Ͻ6�ϽH�ϽB�Ͻy�Ͻ˝Ͻ�ϽŝϽҝϽP   P   ӝϽ��Ͻ͝Ͻ̝Ͻ��Ͻ͝ϽY�Ͻ��Ͻ��Ͻ��Ͻi�Ͻ!�ϽQ�Ͻ7�Ͻ�Ͻ��Ͻy�Ͻ[�Ͻz�ϽR�ϽP   P   �Ͻ�ϽA�Ͻm�ϽH�Ͻ��Ͻ�Ͻ��Ͻ��Ͻc�Ͻi�Ͻ�ϽZ�Ͻ$�Ͻ��Ͻ�ϽB�Ͻ��ϽٝϽ��ϽP   P   -�Ͻ$�ϽR�ϽW�Ͻv�ϽH�Ͻ�Ͻ�Ͻ��ϽҝϽ��Ͻ<�Ͻ<�ϽO�Ͻ$�Ͻ7�ϽH�ϽÝϽ��ϽӝϽP   P   S�Ͻq�Ͻ��Ͻn�Ͻ��ϽP�ϽĞϽ��ϽL�Ͻ��Ͻ��ϽG�Ͻ<�Ͻ<�ϽZ�ϽQ�Ͻ6�ϽN�Ͻ��Ͻ?�ϽP   P   !�ϽM�Ͻ�Ͻ4�ϽD�Ͻ1�ϽW�Ͻ��Ͻ_�ϽK�Ͻ�ϽG�ϽG�Ͻ<�Ͻ�Ͻ!�Ͻ�ϽP�ϽK�Ͻ)�ϽP   P   ��Ͻ��Ͻ��ϽQ�Ͻ̞Ͻ\�Ͻ��Ͻ@�Ͻ�Ͻ��ϽܞϽ�Ͻ��Ͻ��Ͻi�Ͻi�Ͻ:�ϽɝϽ��Ͻ�ϽP   P   v�Ͻs�Ͻ��Ͻ�Ͻ^�ϽI�Ͻm�Ͻ1�Ͻ �Ͻ��Ͻ��ϽK�Ͻ��ϽҝϽc�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   �Ͻm�Ͻ��Ͻ0�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ0�Ͻ �Ͻ�Ͻ_�ϽL�Ͻ��Ͻ��Ͻ��Ͻz�Ͻ��Ͻ|�Ͻ,�ϽP   P   �Ͻ��Ͻ�Ͻ(�Ͻ<�ϽמϽc�Ͻ+�Ͻ�Ͻ1�Ͻ@�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ؝Ͻ-�Ͻ�Ͻ��ϽP   P   ��ϽV�ϽV�Ͻ[�Ͻ��Ͻ�Ͻ��Ͻc�Ͻ��Ͻm�Ͻ��ϽW�ϽĞϽ�Ͻ�ϽY�Ͻ��ϽG�Ͻs�ϽS�ϽP   P   �Ͻ�ϽV�Ͻ��Ͻ`�Ͻ%�Ͻ�ϽמϽ�ϽI�Ͻ\�Ͻ1�ϽP�ϽH�Ͻ��Ͻ͝Ͻ��Ͻ��Ͻk�Ͻ�ϽP   P   ��Ͻ˝Ͻ�Ͻ{�Ͻd�Ͻ`�Ͻ��Ͻ<�Ͻ�Ͻ^�Ͻ̞ϽD�Ͻ��Ͻv�ϽH�Ͻ��Ͻ�Ͻk�Ͻ[�Ͻ��ϽP   P   )�Ͻ�ϽΝϽ��Ͻ{�Ͻ��Ͻ[�Ͻ(�Ͻ0�Ͻ�ϽQ�Ͻ4�Ͻn�ϽW�Ͻm�Ͻ̝Ͻ��Ͻ&�Ͻh�Ͻ��ϽP   P   <�Ͻ}�Ͻ�ϽΝϽ�ϽV�ϽV�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽR�ϽA�Ͻ͝Ͻg�Ͻ^�Ͻp�Ͻ�ϽP   P   a�Ͻ��Ͻ}�Ͻ�Ͻ˝Ͻ�ϽV�Ͻ��Ͻm�Ͻs�Ͻ��ϽM�Ͻq�Ͻ$�Ͻ�Ͻ��Ͻ~�Ͻ��Ͻ�ϽY�ϽP   P   e�Ͻt�Ͻ��Ͻ��ϽX�ϽȟϽ�Ͻ�Ͻ7�ϽG�Ͻ��Ͻ�Ͻk�Ͻ�ϽK�Ͻ��ϽßϽşϽ��Ͻg�ϽP   P   g�ϽR�Ͻk�Ͻ��Ͻ�Ͻ�Ͻ-�Ͻ?�Ͻ	�Ͻ	�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻa�ϽP   P   ��Ͻ��Ͻ��ϽğϽ�Ͻ@�Ͻ��ϽB�Ͻ��Ͻ��Ͻ�Ͻu�Ͻ��Ͻs�Ͻ
�Ͻ(�Ͻ�ϽR�Ͻ�Ͻ��ϽP   P   şϽ��Ͻ��Ͻ��ϽʟϽQ�Ͻ˞ϽO�Ͻ��ϽߟϽ�Ͻ �Ͻ�Ͻ�Ͻ��Ͻ��Ͻ(�Ͻv�ϽR�Ͻ��ϽP   P   ßϽٟϽ�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ�ϽZ�ϽԟϽϽϟϽ�Ͻ՟ϽџϽ��Ͻ��Ͻ(�Ͻ�Ͻ��ϽP   P   ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ;�ϽD�Ͻ͟ϽӟϽ|�Ͻ��ϽşϽşϽ��Ͻ��Ͻ��Ͻ��Ͻ(�Ͻ�ϽP   P   K�Ͻ�Ͻ��Ͻ��Ͻ՟Ͻ6�Ͻ	�Ͻ>�Ͻ��Ͻ��ϽğϽϟϽ��Ͻ��Ͻ��Ͻ��ϽџϽ��Ͻ
�Ͻ�ϽP   P   �Ͻ�ϽF�Ͻ=�Ͻt�Ͻ)�Ͻ,�Ͻ�Ͻ	�Ͻ��Ͻ�ϽݟϽϽ��Ͻ��ϽşϽ՟Ͻ�Ͻs�Ͻ��ϽP   P   k�Ͻ�Ͻy�Ͻ�Ͻ��Ͻ�ϽP�Ͻ �Ͻ.�Ͻ�ϽßϽ�ϽɟϽϽ��ϽşϽ�Ͻ�Ͻ��Ͻ�ϽP   P   �ϽY�Ͻ
�ϽĠϽ��Ͻ~�Ͻ��Ͻ�Ͻa�Ͻ+�Ͻ�Ͻ��Ͻ�ϽݟϽϟϽ��ϽϟϽ �Ͻu�Ͻ��ϽP   P   ��Ͻ,�Ͻ��Ͻ�ϽϠϽu�ϽƠϽ��Ͻn�Ͻ'�Ͻ��Ͻ�ϽßϽ�ϽğϽ|�ϽϽ�Ͻ�Ͻ��ϽP   P   G�Ͻ"�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ)�Ͻ�Ͻ��Ͻ��Ͻ'�Ͻ+�Ͻ�Ͻ��Ͻ��ϽӟϽԟϽߟϽ��Ͻ	�ϽP   P   7�Ͻ0�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��Ͻn�Ͻa�Ͻ.�Ͻ	�Ͻ��Ͻ͟ϽZ�Ͻ��Ͻ��Ͻ	�ϽP   P   �Ͻ/�Ͻ�Ͻ�Ͻ�Ͻ�ϽT�ϽA�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ �Ͻ�Ͻ>�ϽD�Ͻ�ϽO�ϽB�Ͻ?�ϽP   P   �Ͻ1�Ͻ;�ϽʠϽԠϽ$�Ͻ��ϽT�Ͻ�Ͻ)�ϽƠϽ��ϽP�Ͻ,�Ͻ	�Ͻ;�Ͻ��Ͻ˞Ͻ��Ͻ-�ϽP   P   ȟϽB�Ͻ9�Ͻ2�Ͻ��Ͻk�Ͻ$�Ͻ�Ͻ��Ͻ�Ͻu�Ͻ~�Ͻ�Ͻ)�Ͻ6�Ͻ��Ͻ�ϽQ�Ͻ@�Ͻ�ϽP   P   X�Ͻ��Ͻ˟ϽZ�Ͻd�Ͻ��ϽԠϽ�Ͻ�Ͻ�ϽϠϽ��Ͻ��Ͻt�Ͻ՟Ͻ��Ͻ��ϽʟϽ�Ͻ�ϽP   P   ��Ͻ�Ͻ�Ͻ��ϽZ�Ͻ2�ϽʠϽ�Ͻ�Ͻ�Ͻ�ϽĠϽ�Ͻ=�Ͻ��Ͻ�Ͻ�Ͻ��ϽğϽ��ϽP   P   ��Ͻ��ϽǟϽ�Ͻ˟Ͻ9�Ͻ;�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ
�Ͻy�ϽF�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻk�ϽP   P   t�Ͻ^�Ͻ��Ͻ�Ͻ��ϽB�Ͻ1�Ͻ/�Ͻ0�Ͻ"�Ͻ,�ϽY�Ͻ�Ͻ�Ͻ�Ͻ��ϽٟϽ��Ͻ��ϽR�ϽP   P   �ϽޡϽ�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ@�Ͻ'�Ͻw�Ͻ��Ͻh�Ͻ�Ͻ*�Ͻ�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ�ϽP   P   �Ͻ�ϽK�Ͻ8�Ͻ��Ͻ��Ͻ��Ͻ��ϽۡϽ�Ͻ��Ͻ)�ϽڡϽ�Ͻ��Ͻg�Ͻ��Ͻ��Ͻk�Ͻ<�ϽP   P   ��Ͻc�ϽԡϽ��Ͻ��ϽH�Ͻ�Ͻq�Ͻ��ϽS�Ͻ��Ͻ�Ͻ��ϽD�Ͻ�Ͻf�Ͻ5�ϽQ�Ͻ��Ͻk�ϽP   P   ��Ͻ��Ͻ͡Ͻ�Ͻ��Ͻ/�Ͻ͢Ͻ2�Ͻ֡Ͻ�Ͻ{�Ͻj�ϽD�Ͻ��ϽѡϽ�Ͻ0�Ͻ��ϽQ�Ͻ��ϽP   P   �Ͻ¡Ͻ��ϽΡϽ��Ͻ��Ͻ�Ͻ5�Ͻ;�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ~�Ͻ��Ͻ��Ͻ:�Ͻ0�Ͻ5�Ͻ��ϽP   P   �Ͻ?�Ͻ=�Ͻ&�Ͻs�Ͻ�Ͻp�Ͻr�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻf�Ͻg�ϽP   P   �Ͻ�Ͻ8�Ͻ�Ͻ �Ͻ#�ϽáϽ��ϽšϽ�Ͻ��Ͻ��Ͻ�Ͻ=�Ͻ��Ͻ��Ͻ��ϽѡϽ�Ͻ��ϽP   P   *�Ͻ:�Ͻ~�ϽF�Ͻj�Ͻ\�Ͻc�ϽD�Ͻ��Ͻ^�Ͻ��Ͻ��Ͻ��ϽC�Ͻ=�Ͻ��Ͻ~�Ͻ��ϽD�Ͻ�ϽP   P   �Ͻ.�ϽL�Ͻ��Ͻp�Ͻ��Ͻ�Ͻ9�Ͻ�Ͻ�Ͻ��Ͻe�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽD�Ͻ��ϽڡϽP   P   h�ϽY�ϽšϽ��Ͻ��Ͻr�Ͻ��ϽۡϽj�Ͻr�Ͻ �Ͻ��Ͻe�Ͻ��Ͻ��Ͻ��Ͻ��Ͻj�Ͻ�Ͻ)�ϽP   P   ��Ͻ��ϽY�Ͻ��Ͻ�Ͻ��ϽۢϽ��Ͻ/�Ͻ�ϽN�Ͻ �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ{�Ͻ��Ͻ��ϽP   P   w�Ͻ�Ͻ��Ͻc�ϽK�Ͻ��Ͻ}�ϽN�Ͻf�Ͻ��Ͻ�Ͻr�Ͻ�Ͻ^�Ͻ�Ͻ��Ͻ��Ͻ�ϽS�Ͻ�ϽP   P   '�Ͻ5�Ͻj�ϽE�Ͻw�ϽI�ϽˢϽL�Ͻa�Ͻf�Ͻ/�Ͻj�Ͻ�Ͻ��ϽšϽ�Ͻ;�Ͻ֡Ͻ��ϽۡϽP   P   @�Ͻ1�ϽޡϽ��ϽP�ϽK�Ͻ8�Ͻ`�ϽL�ϽN�Ͻ��ϽۡϽ9�ϽD�Ͻ��Ͻr�Ͻ5�Ͻ2�Ͻq�Ͻ��ϽP   P   �Ͻ)�ϽK�Ͻ��Ͻ��ϽZ�Ͻ�Ͻ8�ϽˢϽ}�ϽۢϽ��Ͻ�Ͻc�ϽáϽp�Ͻ�Ͻ͢Ͻ�Ͻ��ϽP   P   ��Ͻ"�Ͻ[�Ͻ��Ͻz�Ͻ¢ϽZ�ϽK�ϽI�Ͻ��Ͻ��Ͻr�Ͻ��Ͻ\�Ͻ#�Ͻ�Ͻ��Ͻ/�ϽH�Ͻ��ϽP   P   �ϽY�Ͻ-�ϽI�Ͻ��Ͻz�Ͻ��ϽP�Ͻw�ϽK�Ͻ�Ͻ��Ͻp�Ͻj�Ͻ �Ͻs�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ0�Ͻ��ϽI�Ͻ��Ͻ��Ͻ��ϽE�Ͻc�Ͻ��Ͻ��Ͻ��ϽF�Ͻ�Ͻ&�ϽΡϽ�Ͻ��Ͻ8�ϽP   P   �Ͻ��Ͻ��Ͻ0�Ͻ-�Ͻ[�ϽK�ϽޡϽj�Ͻ��ϽY�ϽšϽL�Ͻ~�Ͻ8�Ͻ=�Ͻ��Ͻ͡ϽԡϽK�ϽP   P   ޡϽ�Ͻ��Ͻ��ϽY�Ͻ"�Ͻ)�Ͻ1�Ͻ5�Ͻ�Ͻ��ϽY�Ͻ.�Ͻ:�Ͻ�Ͻ?�Ͻ¡Ͻ��Ͻc�Ͻ�ϽP   P   ��ϽݣϽ��ϽޣϽU�Ͻ1�Ͻ1�Ͻj�Ͻ�Ͻ�Ͻ �Ͻ�Ͻ�Ͻ2�Ͻ�Ͻ]�Ͻ��Ͻ�Ͻ�ϽأϽP   P   أϽ�ϽR�Ͻ�Ͻ�Ͻ�Ͻ��ϽK�Ͻ�Ͻ�Ͻ>�Ͻ�Ͻ�Ͻ$�Ͻ��Ͻp�Ͻ�Ͻ<�Ͻ��Ͻm�ϽP   P   �Ͻ
�Ͻ[�Ͻ�Ͻ�Ͻm�ϽڣϽ��Ͻ5�Ͻ�Ͻ�ϽӣϽ�Ͻ�Ͻ�Ͻ�Ͻ��Ͻm�ϽڣϽ��ϽP   P   �ϽK�ϽB�Ͻ�Ͻ�Ͻi�ϽW�Ͻp�Ͻ�Ͻ��Ͻ��ϽM�Ͻ\�Ͻ��ϽˣϽ�Ͻ��ϽY�Ͻm�Ͻ<�ϽP   P   ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ4�Ͻ��Ͻ��ϽΣϽ��ϽT�Ͻb�Ͻi�ϽC�Ͻ'�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   ]�Ͻ�Ͻ�Ͻ��ϽݣϽe�ϽT�Ͻ.�Ͻ�ϽϣϽZ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ'�Ͻ�Ͻ�Ͻ�Ͻp�ϽP   P   �Ͻ��Ͻ�Ͻm�Ͻ�Ͻ��Ͻ�Ͻs�Ͻ�ϽУϽ(�ϽɣϽ��Ͻ�Ͻg�Ͻ�Ͻ'�ϽˣϽ�Ͻ��ϽP   P   2�Ͻ�Ͻ	�Ͻ%�Ͻ�Ͻ�Ͻ�ϽO�Ͻ�Ͻ�Ͻ
�Ͻ;�Ͻ��Ͻ��Ͻ�Ͻ��ϽC�Ͻ��Ͻ�Ͻ$�ϽP   P   �Ͻ�ϽQ�ϽM�Ͻ�Ͻf�Ͻg�Ͻ��Ͻ
�Ͻ�Ͻ�ϽR�Ͻq�Ͻ��Ͻ��Ͻ��Ͻi�Ͻ\�Ͻ�Ͻ�ϽP   P   �Ͻ��Ͻ\�Ͻ�ϽM�ϽV�Ͻ��Ͻ��Ͻw�Ͻ�Ͻ*�Ͻ�ϽR�Ͻ;�ϽɣϽ��Ͻb�ϽM�ϽӣϽ�ϽP   P    �Ͻ��Ͻ��Ͻ��Ͻ:�Ͻ��Ͻ^�Ͻ��Ͻ��Ͻ��Ͻ
�Ͻ*�Ͻ�Ͻ
�Ͻ(�ϽZ�ϽT�Ͻ��Ͻ�Ͻ>�ϽP   P   �Ͻ��Ͻ	�Ͻ�Ͻ��Ͻ�ϽʤϽ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�Ͻ�ϽУϽϣϽ��Ͻ��Ͻ�Ͻ�ϽP   P   �Ͻ��Ͻ��Ͻ�ϽפϽa�Ͻ6�ϽE�Ͻ��Ͻ��Ͻ��Ͻw�Ͻ
�Ͻ�Ͻ�Ͻ�ϽΣϽ�Ͻ5�Ͻ�ϽP   P   j�Ͻ��Ͻp�Ͻ��Ͻ��Ͻ8�Ͻ~�Ͻ��ϽE�Ͻ��Ͻ��Ͻ��Ͻ��ϽO�Ͻs�Ͻ.�Ͻ��Ͻp�Ͻ��ϽK�ϽP   P   1�Ͻ�Ͻ��Ͻ��Ͻd�ϽƤϽ��Ͻ~�Ͻ6�ϽʤϽ^�Ͻ��Ͻg�Ͻ�Ͻ�ϽT�Ͻ��ϽW�ϽڣϽ��ϽP   P   1�Ͻ��Ͻ�Ͻ>�Ͻ=�Ͻ�ϽƤϽ8�Ͻa�Ͻ�Ͻ��ϽV�Ͻf�Ͻ�Ͻ��Ͻe�Ͻ4�Ͻi�Ͻm�Ͻ�ϽP   P   U�ϽݣϽ$�Ͻ�ϽR�Ͻ=�Ͻd�Ͻ��ϽפϽ��Ͻ:�ϽM�Ͻ�Ͻ�Ͻ�ϽݣϽ�Ͻ�Ͻ�Ͻ�ϽP   P   ޣϽe�ϽأϽl�Ͻ�Ͻ>�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�ϽM�Ͻ%�Ͻm�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�ϽP   P   ��Ͻ8�Ͻ1�ϽأϽ$�Ͻ�Ͻ��Ͻp�Ͻ��Ͻ	�Ͻ��Ͻ\�ϽQ�Ͻ	�Ͻ�Ͻ�Ͻ�ϽB�Ͻ[�ϽR�ϽP   P   ݣϽ�Ͻ8�Ͻe�ϽݣϽ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻ��ϽK�Ͻ
�Ͻ�ϽP   P   ��ϽԥϽ�ϽԥϽ�Ͻ��Ͻ	�Ͻ֥ϽC�ϽF�Ͻq�Ͻq�Ͻ	�Ͻ��ϽեϽ��Ͻ��ϽɥϽեϽץϽP   P   ץϽ�Ͻ�ϽX�Ͻ��ϽĥϽ�Ͻ��Ͻ'�ϽE�ϽO�Ͻ
�Ͻp�ϽC�Ͻ�ϽإϽ��Ͻ�ϽD�Ͻ>�ϽP   P   եϽ��Ͻ�ϽI�Ͻ
�ϽG�Ͻp�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ	�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�ϽJ�Ͻ˥ϽD�ϽP   P   ɥϽ٥Ͻ��Ͻ��Ͻ��ϽB�ϽD�Ͻ�Ͻk�ϽѥϽ��Ͻ��Ͻ�ϽۥϽ�ϽU�Ͻ?�Ͻ��ϽJ�Ͻ�ϽP   P   ��Ͻe�ϽH�ϽV�Ͻ�Ͻ�ϽU�Ͻ3�Ͻ�Ͻ�Ͻ�Ͻ��ϽG�Ͻ��Ͻ��Ͻ!�Ͻ��Ͻ?�Ͻ�Ͻ��ϽP   P   ��ϽG�Ͻ��Ͻ/�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�ϽΥϽ��ϽA�Ͻ%�Ͻ"�Ͻ��Ͻ!�ϽU�Ͻ�ϽإϽP   P   եϽ��Ͻ5�Ͻ�ϽV�Ͻ��Ͻ,�Ͻ٥Ͻ��Ͻ�ϽʥϽ��Ͻ��Ͻ��Ͻ=�Ͻ"�Ͻ��Ͻ�Ͻ��Ͻ�ϽP   P   ��ϽQ�Ͻ]�Ͻc�Ͻ�Ͻy�Ͻ$�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��ϽM�Ͻ<�Ͻ��Ͻ%�Ͻ��ϽۥϽ�ϽC�ϽP   P   	�Ͻ�Ͻ�Ͻo�Ͻz�ϽX�ϽB�Ͻ��Ͻz�Ͻ^�Ͻ'�ϽХϽ^�ϽM�Ͻ��ϽA�ϽG�Ͻ�Ͻ��Ͻp�ϽP   P   q�Ͻ�ϽD�ϽߦϽ��ϽæϽ��Ͻ~�Ͻ�Ͻ9�Ͻ�Ͻ��ϽХϽ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ	�Ͻ
�ϽP   P   q�Ͻ��ϽQ�Ͻ��Ͻ)�Ͻ�Ͻ?�ϽL�Ͻj�Ͻ��ϽæϽ�Ͻ'�Ͻ�ϽʥϽΥϽ�Ͻ��Ͻ��ϽO�ϽP   P   F�Ͻ��Ͻ��Ͻ�Ͻ~�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ9�Ͻ^�Ͻ��Ͻ�Ͻ�Ͻ�ϽѥϽ�ϽE�ϽP   P   C�Ͻ<�ϽT�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ|�Ͻ�Ͻj�Ͻ�Ͻz�Ͻ�Ͻ��Ͻ�Ͻ�Ͻk�Ͻ��Ͻ'�ϽP   P   ֥Ͻ��Ͻf�Ͻ\�Ͻ��Ͻi�Ͻ��ϽզϽ��Ͻ��ϽL�Ͻ~�Ͻ��Ͻ��Ͻ٥Ͻ�Ͻ3�Ͻ�Ͻ�Ͻ��ϽP   P   	�Ͻ"�ϽT�ϽѦϽ@�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ?�Ͻ��ϽB�Ͻ$�Ͻ,�Ͻ��ϽU�ϽD�Ͻp�Ͻ�ϽP   P   ��Ͻ��Ͻg�Ͻ3�Ͻ��Ͻ�Ͻ��Ͻi�Ͻ��Ͻ��Ͻ�ϽæϽX�Ͻy�Ͻ��Ͻ��Ͻ�ϽB�ϽG�ϽĥϽP   P   �Ͻ-�ϽX�Ͻ3�Ͻ��Ͻ��Ͻ@�Ͻ��Ͻ��Ͻ~�Ͻ)�Ͻ��Ͻz�Ͻ�ϽV�Ͻ�Ͻ�Ͻ��Ͻ
�Ͻ��ϽP   P   ԥϽ;�Ͻ
�Ͻ%�Ͻ3�Ͻ3�ϽѦϽ\�Ͻ�Ͻ�Ͻ��ϽߦϽo�Ͻc�Ͻ�Ͻ/�ϽV�Ͻ��ϽI�ϽX�ϽP   P   �Ͻ��Ͻ��Ͻ
�ϽX�Ͻg�ϽT�Ͻf�ϽT�Ͻ��ϽQ�ϽD�Ͻ�Ͻ]�Ͻ5�Ͻ��ϽH�Ͻ��Ͻ�Ͻ�ϽP   P   ԥϽ�Ͻ��Ͻ;�Ͻ-�Ͻ��Ͻ"�Ͻ��Ͻ<�Ͻ��Ͻ��Ͻ�Ͻ�ϽQ�Ͻ��ϽG�Ͻe�Ͻ٥Ͻ��Ͻ�ϽP   P   *�Ͻ�Ͻb�Ͻ6�Ͻ_�Ͻ�Ͻd�Ͻ~�Ͻ��Ͻ�Ͻ�Ͻ�Ͻq�Ͻt�ϽH�Ͻ�Ͻ4�Ͻ+�ϽU�Ͻ�ϽP   P   �Ͻ�Ͻ��Ͻ��ϽاϽG�Ͻ/�ϽE�ϽN�Ͻ�Ͻ�Ͻ�Ͻ�Ͻ]�Ͻ`�Ͻ4�Ͻd�Ͻ��Ͻ��Ͻ�ϽP   P   U�Ͻ�Ͻj�Ͻ��Ͻ��ϽD�Ͻ�ϽçϽ/�ϽH�Ͻ�ϽX�Ͻ��ϽN�Ͻ�Ͻ�Ͻ��Ͻ �Ͻ��Ͻ��ϽP   P   +�Ͻ�ϽƧϽ�Ͻ�Ͻ#�Ͻ��Ͻ�Ͻ�Ͻ:�Ͻ`�Ͻ4�ϽN�ϽK�ϽQ�Ͻ��Ͻ�Ͻ�Ͻ �Ͻ��ϽP   P   4�ϽA�Ͻ��Ͻ=�ϽW�ϽZ�Ͻ�Ͻ.�Ͻ�Ͻ��Ͻ-�Ͻ7�Ͻ)�Ͻ2�Ͻ�Ͻ�ϽӧϽ�Ͻ��Ͻd�ϽP   P   �Ͻ�Ͻ �Ͻ�Ͻ�Ͻ�Ͻ�ϽЧϽħϽ�Ͻ4�ϽէϽ,�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻ4�ϽP   P   H�Ͻ&�ϽɧϽ#�ϽߧϽ�Ͻ��ϽI�ϽN�Ͻg�Ͻ�Ͻ�Ͻ�ϽC�Ͻ�Ͻ��Ͻ�ϽQ�Ͻ�Ͻ`�ϽP   P   t�Ͻr�Ͻ�Ͻr�Ͻ^�Ͻ�ϽY�ϽX�Ͻ=�Ͻ%�ϽK�ϽA�Ͻ#�Ͻ�ϽC�Ͻ�Ͻ2�ϽK�ϽN�Ͻ]�ϽP   P   q�Ͻ��Ͻ�Ͻ��Ͻ �Ͻ�Ͻ4�Ͻ|�Ͻ��Ͻ�Ͻ8�ϽL�Ͻ�Ͻ#�Ͻ�Ͻ,�Ͻ)�ϽN�Ͻ��Ͻ�ϽP   P   �ϽC�Ͻ+�Ͻ]�Ͻ.�Ͻl�ϽO�Ͻ@�Ͻ0�ϽߧϽ�Ͻ5�ϽL�ϽA�Ͻ�ϽէϽ7�Ͻ4�ϽX�Ͻ�ϽP   P   �Ͻ�Ͻ0�ϽH�Ͻ��Ͻv�Ͻ��Ͻ1�Ͻ>�Ͻ�Ͻ�Ͻ�Ͻ8�ϽK�Ͻ�Ͻ4�Ͻ-�Ͻ`�Ͻ�Ͻ�ϽP   P   �Ͻ�Ͻ��Ͻf�Ͻb�ϽU�Ͻ6�Ͻ��Ͻc�Ͻ��Ͻ�ϽߧϽ�Ͻ%�Ͻg�Ͻ�Ͻ��Ͻ:�ϽH�Ͻ�ϽP   P   ��Ͻ<�Ͻ!�Ͻ]�Ͻ��Ͻo�ϽZ�Ͻ`�ϽY�Ͻc�Ͻ>�Ͻ0�Ͻ��Ͻ=�ϽN�ϽħϽ�Ͻ�Ͻ/�ϽN�ϽP   P   ~�Ͻ|�Ͻ2�Ͻ;�Ͻm�Ͻc�Ͻj�Ͻu�Ͻ`�Ͻ��Ͻ1�Ͻ@�Ͻ|�ϽX�ϽI�ϽЧϽ.�Ͻ�ϽçϽE�ϽP   P   d�Ͻe�Ͻ7�ϽO�Ͻ��ϽF�Ͻp�Ͻj�ϽZ�Ͻ6�Ͻ��ϽO�Ͻ4�ϽY�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻ/�ϽP   P   �Ͻ�Ͻ�Ͻ�ϽJ�Ͻv�ϽF�Ͻc�Ͻo�ϽU�Ͻv�Ͻl�Ͻ�Ͻ�Ͻ�Ͻ�ϽZ�Ͻ#�ϽD�ϽG�ϽP   P   _�Ͻ�Ͻ֧Ͻ_�Ͻ#�ϽJ�Ͻ��Ͻm�Ͻ��Ͻb�Ͻ��Ͻ.�Ͻ �Ͻ^�ϽߧϽ�ϽW�Ͻ�Ͻ��ϽاϽP   P   6�Ͻ$�Ͻ�Ͻ+�Ͻ_�Ͻ�ϽO�Ͻ;�Ͻ]�Ͻf�ϽH�Ͻ]�Ͻ��Ͻr�Ͻ#�Ͻ�Ͻ=�Ͻ�Ͻ��Ͻ��ϽP   P   b�ϽƧϽݧϽ�Ͻ֧Ͻ�Ͻ7�Ͻ2�Ͻ!�Ͻ��Ͻ0�Ͻ+�Ͻ�Ͻ�ϽɧϽ �Ͻ��ϽƧϽj�Ͻ��ϽP   P   �Ͻ1�ϽƧϽ$�Ͻ�Ͻ�Ͻe�Ͻ|�Ͻ<�Ͻ�Ͻ�ϽC�Ͻ��Ͻr�Ͻ&�Ͻ�ϽA�Ͻ�Ͻ�Ͻ�ϽP   P   ��ϽݩϽ�Ͻ�ϽکϽR�Ͻ�Ͻ��ϽթϽ��Ͻ��Ͻr�Ͻ�ϽީϽ��Ͻ7�Ͻ�Ͻ�Ͻ��Ͻ۩ϽP   P   ۩Ͻ��Ͻ�ϽI�ϽI�Ͻ��ϽN�ϽA�Ͻ©Ͻ2�ϽO�Ͻ��Ͻ�Ͻ��Ͻ
�ϽX�Ͻ�Ͻ"�Ͻ\�Ͻ��ϽP   P   ��ϽܩϽ�Ͻg�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ*�Ͻ
�Ͻ0�Ͻ5�ϽB�Ͻi�Ͻ�Ͻ�Ͻ �Ͻ\�ϽP   P   �Ͻf�Ͻ��Ͻ�Ͻo�ϽҩϽʩϽd�Ͻ�Ͻ��Ͻ��Ͻ�ϽƩϽ٩Ͻ��Ͻ�ϽG�Ͻ�Ͻ�Ͻ"�ϽP   P   �Ͻ��ϽI�ϽթϽ�Ͻ
�Ͻ �Ͻu�Ͻ�Ͻ&�ϽҩϽ9�Ͻm�ϽQ�Ͻ��Ͻ	�Ͻ:�ϽG�Ͻ�Ͻ�ϽP   P   7�Ͻ�Ͻ��Ͻ\�ϽO�Ͻ3�Ͻo�ϽP�Ͻ��Ͻ(�ϽV�Ͻj�Ͻ��Ͻ��Ͻ"�Ͻ}�Ͻ	�Ͻ�Ͻi�ϽX�ϽP   P   ��Ͻ��Ͻp�Ͻ?�ϽN�Ͻ�Ͻ�Ͻ6�Ͻ-�Ͻ�ϽΩϽA�Ͻ�Ͻ!�Ͻ��Ͻ"�Ͻ��Ͻ��ϽB�Ͻ
�ϽP   P   ީϽ�Ͻf�ϽC�Ͻo�Ͻ]�Ͻ��Ͻ̩ϽөϽ�Ͻ��Ͻl�Ͻ��Ͻj�Ͻ!�Ͻ��ϽQ�Ͻ٩Ͻ5�Ͻ��ϽP   P   �Ͻ�Ͻ��Ͻ��ϽY�Ͻ��Ͻv�ϽP�ϽЩϽ/�Ͻ%�Ͻ��Ͻ3�Ͻ��Ͻ�Ͻ��Ͻm�ϽƩϽ0�Ͻ�ϽP   P   r�Ͻ~�Ͻm�Ͻ
�Ͻ+�Ͻ?�Ͻ/�ϽK�Ͻ��Ͻq�Ͻ��ϽީϽ��Ͻl�ϽA�Ͻj�Ͻ9�Ͻ�Ͻ
�Ͻ��ϽP   P   ��Ͻ�Ͻ~�ϽU�Ͻn�ϽΪϽ@�Ͻv�Ͻl�Ͻ�Ͻp�Ͻ��Ͻ%�Ͻ��ϽΩϽV�ϽҩϽ��Ͻ*�ϽO�ϽP   P   ��Ͻ�Ͻ �Ͻ��ϽI�ϽY�Ͻl�ϽX�Ͻ��Ͻ�Ͻ�Ͻq�Ͻ/�Ͻ�Ͻ�Ͻ(�Ͻ&�Ͻ��Ͻ�Ͻ2�ϽP   P   թϽI�Ͻ��Ͻ��ϽX�ϽQ�Ͻ��Ͻr�ϽE�Ͻ��Ͻl�Ͻ��ϽЩϽөϽ-�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ©ϽP   P   ��Ͻe�Ͻj�Ͻ��Ͻ>�Ͻ��ϽY�ϽF�Ͻr�ϽX�Ͻv�ϽK�ϽP�Ͻ̩Ͻ6�ϽP�Ͻu�Ͻd�Ͻ�ϽA�ϽP   P   �Ͻ�Ͻf�Ͻ��Ͻb�Ͻe�Ͻk�ϽY�Ͻ��Ͻl�Ͻ@�Ͻ/�Ͻv�Ͻ��Ͻ�Ͻo�Ͻ �ϽʩϽ��ϽN�ϽP   P   R�Ͻ�Ͻf�ϽͪϽ2�ϽͪϽe�Ͻ��ϽQ�ϽY�ϽΪϽ?�Ͻ��Ͻ]�Ͻ�Ͻ3�Ͻ
�ϽҩϽ�Ͻ��ϽP   P   کϽ>�Ͻ\�ϽM�Ͻ5�Ͻ2�Ͻb�Ͻ>�ϽX�ϽI�Ͻn�Ͻ+�ϽY�Ͻo�ϽN�ϽO�Ͻ�Ͻo�Ͻ��ϽI�ϽP   P   �Ͻ��Ͻ��ϽS�ϽM�ϽͪϽ��Ͻ��Ͻ��Ͻ��ϽU�Ͻ
�Ͻ��ϽC�Ͻ?�Ͻ\�ϽթϽ�Ͻg�ϽI�ϽP   P   �Ͻ��ϽG�Ͻ��Ͻ\�Ͻf�Ͻf�Ͻj�Ͻ��Ͻ �Ͻ~�Ͻm�Ͻ��Ͻf�Ͻp�Ͻ��ϽI�Ͻ��Ͻ�Ͻ�ϽP   P   ݩϽ��Ͻ��Ͻ��Ͻ>�Ͻ�Ͻ�Ͻe�ϽI�Ͻ�Ͻ�Ͻ~�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ��Ͻf�ϽܩϽ��ϽP   P   ��Ͻ{�Ͻ�Ͻ-�Ͻ5�ϽI�ϽS�Ͻ��ϽB�ϽH�Ͻ�Ͻ�Ͻ}�Ͻ�Ͻy�Ͻ �Ͻ��Ͻ.�Ͻ+�Ͻ��ϽP   P   ��Ͻe�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��Ͻ#�Ͻ��Ͻ��Ͻ��ϽϫϽ]�Ͻ��Ͻ�ϽϫϽ��Ͻ��Ͻ�Ͻy�ϽP   P   +�Ͻ�Ͻ��ϽޫϽ��ϽJ�Ͻb�Ͻ�Ͻ��Ͻ"�Ͻd�ϽE�Ͻg�Ͻ=�ϽG�Ͻ��Ͻ��Ͻ2�Ͻ�Ͻ�ϽP   P   .�Ͻ�Ͻ%�Ͻ�Ͻ�ϽD�ϽլϽ��Ͻ�Ͻ��Ͻ]�ϽB�Ͻ�Ͻ]�Ͻ]�Ͻ-�Ͻ׫ϽɬϽ2�Ͻ��ϽP   P   ��Ͻ�Ͻ'�Ͻ�Ͻ9�Ͻ�Ͻd�Ͻ�Ͻ��Ͻj�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ&�Ͻ=�ϽH�Ͻ׫Ͻ��Ͻ��ϽP   P    �Ͻ�Ͻ�ϽثϽr�Ͻ/�Ͻ�Ͻ�ϽL�Ͻb�Ͻw�Ͻ�ϽY�Ͻ^�Ͻ�Ͻ��Ͻ=�Ͻ-�Ͻ��ϽϫϽP   P   y�Ͻ��Ͻi�ϽϫϽP�Ͻ��Ͻ6�Ͻ
�Ͻ��Ͻ|�Ͻ�Ͻ<�Ͻd�Ͻ%�ϽάϽ�Ͻ&�Ͻ]�ϽG�Ͻ�ϽP   P   �Ͻa�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��ϽϬϽ��ϽU�ϽL�Ͻ �ϽG�Ͻ��Ͻ%�Ͻ^�Ͻ�Ͻ]�Ͻ=�Ͻ��ϽP   P   }�Ͻ�Ͻ-�ϽR�Ͻb�Ͻ<�Ͻ�Ͻ�Ͻ1�Ͻm�ϽN�Ͻ3�ϽݫϽG�Ͻd�ϽY�Ͻ��Ͻ�Ͻg�Ͻ]�ϽP   P   �Ͻ�Ͻ9�Ͻ:�ϽK�Ͻ8�Ͻy�Ͻ��Ͻ%�Ͻ=�ϽǫϽ8�Ͻ3�Ͻ �Ͻ<�Ͻ�Ͻ�ϽB�ϽE�ϽϫϽP   P   �Ͻ��ϽD�Ͻ;�Ͻ`�Ͻ�Ͻ5�Ͻ`�Ͻ<�Ͻ��Ͻ׫ϽǫϽN�ϽL�Ͻ�Ͻw�Ͻ�Ͻ]�Ͻd�Ͻ��ϽP   P   H�Ͻ��Ͻ*�Ͻ�Ͻk�Ͻ�ϽA�Ͻ3�Ͻ�Ͻ&�Ͻ��Ͻ=�Ͻm�ϽU�Ͻ|�Ͻb�Ͻj�Ͻ��Ͻ"�Ͻ��ϽP   P   B�Ͻ�Ͻ@�Ͻ�Ͻ7�Ͻv�Ͻ��Ͻ��Ͻ8�Ͻ�Ͻ<�Ͻ%�Ͻ1�Ͻ��Ͻ��ϽL�Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ��ϽH�Ͻ$�Ͻ[�ϽB�Ͻ��Ͻr�Ͻ0�Ͻ��Ͻ3�Ͻ`�Ͻ��Ͻ�ϽϬϽ
�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ#�ϽP   P   S�Ͻ��Ͻ֫ϽK�Ͻ9�Ͻ?�Ͻe�Ͻr�Ͻ��ϽA�Ͻ5�Ͻy�Ͻ�Ͻ��Ͻ6�Ͻ�Ͻd�ϽլϽb�Ͻ��ϽP   P   I�Ͻ��Ͻ�Ͻ��Ͻ[�Ͻ �Ͻ?�Ͻ��Ͻv�Ͻ�Ͻ�Ͻ8�Ͻ<�Ͻ�Ͻ��Ͻ/�Ͻ�ϽD�ϽJ�Ͻ�ϽP   P   5�ϽJ�ϽE�Ͻ׫Ͻ�Ͻ[�Ͻ9�ϽB�Ͻ7�Ͻk�Ͻ`�ϽK�Ͻb�Ͻ�ϽP�Ͻr�Ͻ9�Ͻ�Ͻ��Ͻ�ϽP   P   -�Ͻ+�Ͻ��ϽȫϽ׫Ͻ��ϽK�Ͻ[�Ͻ�Ͻ�Ͻ;�Ͻ:�ϽR�Ͻ��ϽϫϽثϽ�Ͻ�ϽޫϽ�ϽP   P   �Ͻ�Ͻ�Ͻ��ϽE�Ͻ�Ͻ֫Ͻ$�Ͻ@�Ͻ*�ϽD�Ͻ9�Ͻ-�Ͻ�Ͻi�Ͻ�Ͻ'�Ͻ%�Ͻ��Ͻ��ϽP   P   {�Ͻ�Ͻ�Ͻ+�ϽJ�Ͻ��Ͻ��ϽH�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ�Ͻa�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ�Ͻe�ϽP   P   :�Ͻ�Ͻ�Ͻ]�Ͻ(�Ͻ-�Ͻ"�Ͻ­Ͻ��Ͻ3�Ͻ+�Ͻ-�Ͻ<�Ͻ�Ͻ&�Ͻ�Ͻ~�Ͻc�Ͻ*�Ͻ�ϽP   P   �Ͻ%�Ͻ�Ͻw�Ͻg�Ͻ��Ͻl�Ͻ@�Ͻ?�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ*�Ͻv�Ͻc�ϽP�ϽA�ϽۭϽP   P   *�Ͻ^�Ͻ�Ͻ7�Ͻ*�Ͻ��Ͻ��Ͻ�Ͻ!�Ͻ��Ͻ�Ͻ|�Ͻ �Ͻ��ϽO�Ͻe�Ͻ�Ͻ�Ͻp�ϽA�ϽP   P   c�Ͻ��Ͻ�Ͻ��Ͻm�ϽA�Ͻ��Ͻ�Ͻ+�Ͻ'�Ͻx�ϽX�Ͻ]�ϽI�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ�ϽP�ϽP   P   ~�Ͻv�Ͻw�Ͻb�ϽV�ϽI�Ͻ �Ͻ�ϽO�Ͻ�Ͻa�Ͻ�Ͻ=�Ͻ	�Ͻ��Ͻ�Ͻz�Ͻ��Ͻ�Ͻc�ϽP   P   �Ͻ��Ͻ8�Ͻ3�ϽȭϽ,�Ͻ��Ͻ��ϽJ�Ͻ��ϽL�Ͻ'�ϽL�Ͻ)�Ͻ�Ͻ_�Ͻ�Ͻ�Ͻe�Ͻv�ϽP   P   &�Ͻ��Ͻ]�ϽӮϽG�Ͻ٭Ͻ�Ͻ$�Ͻ!�Ͻ�Ͻ��Ͻ��ϽĭϽ��Ͻ�Ͻ�Ͻ��Ͻ�ϽO�Ͻ*�ϽP   P   �Ͻ�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ'�Ͻ��Ͻ�ϽɭϽH�Ͻ��Ͻ.�ϽѭϽ��Ͻ)�Ͻ	�ϽI�Ͻ��Ͻ�ϽP   P   <�Ͻa�Ͻi�Ͻ�Ͻ}�Ͻ	�Ͻc�Ͻ^�Ͻ)�Ͻ�Ͻ��ϽK�ϽV�Ͻ.�ϽĭϽL�Ͻ=�Ͻ]�Ͻ �Ͻ�ϽP   P   -�Ͻ5�Ͻ��ϽI�ϽN�Ͻ6�Ͻm�Ͻ��ϽM�Ͻ?�Ͻ��Ͻ��ϽK�Ͻ��Ͻ��Ͻ'�Ͻ�ϽX�Ͻ|�Ͻ��ϽP   P   +�Ͻ �Ͻ:�Ͻ5�Ͻ��Ͻ��Ͻ��ϽB�Ͻ;�Ͻ��Ͻ4�Ͻ��Ͻ��ϽH�Ͻ��ϽL�Ͻa�Ͻx�Ͻ�Ͻ��ϽP   P   3�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ@�Ͻz�Ͻk�Ͻ��Ͻ��Ͻ��Ͻ?�Ͻ�ϽɭϽ�Ͻ��Ͻ�Ͻ'�Ͻ��Ͻ�ϽP   P   ��ϽY�Ͻ(�Ͻ��Ͻ��Ͻ�Ͻ@�Ͻ)�Ͻ��Ͻ��Ͻ;�ϽM�Ͻ)�Ͻ�Ͻ!�ϽJ�ϽO�Ͻ+�Ͻ!�Ͻ?�ϽP   P   ­Ͻ��Ͻ��Ͻ5�Ͻ��Ͻ
�ϽP�Ͻ	�Ͻ)�Ͻk�ϽB�Ͻ��Ͻ^�Ͻ��Ͻ$�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ@�ϽP   P   "�ϽO�Ͻ�Ͻ|�Ͻn�Ͻ��Ͻ�ϽP�Ͻ@�Ͻz�Ͻ��Ͻm�Ͻc�Ͻ'�Ͻ�Ͻ��Ͻ �Ͻ��Ͻ��Ͻl�ϽP   P   -�Ͻ�Ͻ�Ͻ&�Ͻ]�Ͻf�Ͻ��Ͻ
�Ͻ�Ͻ@�Ͻ��Ͻ6�Ͻ	�Ͻ�Ͻ٭Ͻ,�ϽI�ϽA�Ͻ��Ͻ��ϽP   P   (�Ͻ��ϽF�Ͻ׮Ͻ�Ͻ]�Ͻn�Ͻ��Ͻ��Ͻ��Ͻ��ϽN�Ͻ}�Ͻ��ϽG�ϽȭϽV�Ͻm�Ͻ*�Ͻg�ϽP   P   ]�Ͻ��ϽK�Ͻ��Ͻ׮Ͻ&�Ͻ|�Ͻ5�Ͻ��Ͻ��Ͻ5�ϽI�Ͻ�Ͻ��ϽӮϽ3�Ͻb�Ͻ��Ͻ7�Ͻw�ϽP   P   �Ͻ �Ͻ*�ϽK�ϽF�Ͻ�Ͻ�Ͻ��Ͻ(�Ͻ��Ͻ:�Ͻ��Ͻi�Ͻ�Ͻ]�Ͻ8�Ͻw�Ͻ�Ͻ�Ͻ�ϽP   P   �Ͻ��Ͻ �Ͻ��Ͻ��Ͻ�ϽO�Ͻ��ϽY�Ͻ��Ͻ �Ͻ5�Ͻa�Ͻ�Ͻ��Ͻ��Ͻv�Ͻ��Ͻ^�Ͻ%�ϽP   P   i�Ͻ:�Ͻ*�ϽկϽ��Ͻl�ϽN�Ͻ��ϽJ�ϽZ�Ͻd�Ͻm�ϽE�Ͻ�ϽK�Ͻ`�Ͻ��ϽȯϽP�ϽG�ϽP   P   G�Ͻj�Ͻ�Ͻ��Ͻ�Ͻ5�Ͻ"�Ͻ%�Ͻ��Ͻd�Ͻ��Ͻ<�Ͻ��Ͻ_�ϽK�Ͻ2�Ͻ�Ͻ�ϽY�Ͻ�ϽP   P   P�Ͻ5�ϽG�ϽG�ϽY�ϽH�Ͻ�Ͻ!�Ͻ{�Ͻ��Ͻ,�Ͻ��Ͻ.�ϽǰϽ{�Ͻ�Ͻ�Ͻ[�ϽA�ϽY�ϽP   P   ȯϽG�Ͻ/�Ͻ��ϽۯϽ{�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ\�Ͻ�Ͻ+�Ͻ�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ[�Ͻ�ϽP   P   ��Ͻ#�Ͻ-�Ͻ�ϽۯϽ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻa�Ͻ�Ͻ'�Ͻ��Ͻr�Ͻ��Ͻ�Ͻ�ϽP   P   `�Ͻ��Ͻ�ϽS�Ͻ��Ͻo�Ͻ#�Ͻ*�Ͻ%�Ͻ�Ͻ��Ͻ*�ϽN�Ͻ2�ϽL�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ2�ϽP   P   K�Ͻ��Ͻ&�Ͻ��ϽC�Ͻq�Ͻd�Ͻ�Ͻ��Ͻ��Ͻ;�Ͻ9�Ͻf�Ͻ�Ͻj�ϽL�Ͻ'�Ͻ�Ͻ{�ϽK�ϽP   P   �ϽV�Ͻ��Ͻ�Ͻ��Ͻ��ϽP�Ͻ
�Ͻk�ϽͰϽD�Ͻ��Ͻ<�ϽڰϽ�Ͻ2�Ͻ�Ͻ�ϽǰϽ_�ϽP   P   E�ϽB�ϽS�Ͻb�Ͻ�Ͻt�ϽW�Ͻ�Ͻe�Ͻ]�Ͻ9�Ͻ��Ͻ��Ͻ<�Ͻf�ϽN�Ͻa�Ͻ+�Ͻ.�Ͻ��ϽP   P   m�ϽM�Ͻ�Ͻ�ϽH�Ͻ>�Ͻ��Ͻ3�Ͻb�Ͻi�ϽC�Ͻ��Ͻ��Ͻ��Ͻ9�Ͻ*�Ͻ��Ͻ�Ͻ��Ͻ<�ϽP   P   d�ϽJ�Ͻ@�Ͻ�Ͻ�Ͻ:�Ͻ)�Ͻ�ϽF�Ͻ-�Ͻ��ϽC�Ͻ9�ϽD�Ͻ;�Ͻ��Ͻ�Ͻ\�Ͻ,�Ͻ��ϽP   P   Z�Ͻ(�Ͻ?�Ͻ��Ͻ)�Ͻ>�ϽG�Ͻ
�Ͻ�ϽV�Ͻ-�Ͻi�Ͻ]�ϽͰϽ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻd�ϽP   P   J�Ͻ��Ͻ)�Ͻ*�Ͻ�Ͻ{�Ͻ��Ͻj�Ͻ!�Ͻ�ϽF�Ͻb�Ͻe�Ͻk�Ͻ��Ͻ%�Ͻ��Ͻ�Ͻ{�Ͻ��ϽP   P   ��Ͻ�Ͻ�Ͻ�Ͻ*�ϽK�Ͻ��Ͻ��Ͻj�Ͻ
�Ͻ�Ͻ3�Ͻ�Ͻ
�Ͻ�Ͻ*�Ͻ��Ͻ��Ͻ!�Ͻ%�ϽP   P   N�Ͻk�ϽR�ϽC�Ͻ��ϽT�Ͻ|�Ͻ��Ͻ��ϽG�Ͻ)�Ͻ��ϽW�ϽP�Ͻd�Ͻ#�Ͻ�Ͻ��Ͻ�Ͻ"�ϽP   P   l�Ͻl�Ͻ��ϽI�ϽZ�Ͻ7�ϽT�ϽK�Ͻ{�Ͻ>�Ͻ:�Ͻ>�Ͻt�Ͻ��Ͻq�Ͻo�Ͻ�Ͻ{�ϽH�Ͻ5�ϽP   P   ��Ͻ��Ͻ:�Ͻ��Ͻ�ϽZ�Ͻ��Ͻ*�Ͻ�Ͻ)�Ͻ�ϽH�Ͻ�Ͻ��ϽC�Ͻ��ϽۯϽۯϽX�Ͻ�ϽP   P   կϽM�Ͻ@�Ͻ�Ͻ��ϽI�ϽC�Ͻ�Ͻ*�Ͻ��Ͻ�Ͻ�Ͻb�Ͻ�Ͻ��ϽS�Ͻ�Ͻ��ϽG�Ͻ��ϽP   P   *�Ͻ2�Ͻ��Ͻ@�Ͻ:�Ͻ��ϽR�Ͻ�Ͻ)�Ͻ?�Ͻ@�Ͻ�ϽS�Ͻ��Ͻ&�Ͻ�Ͻ-�Ͻ/�ϽG�Ͻ�ϽP   P   :�Ͻo�Ͻ2�ϽM�Ͻ��Ͻl�Ͻk�Ͻ�Ͻ��Ͻ(�ϽJ�ϽM�ϽB�ϽV�Ͻ��Ͻ��Ͻ#�ϽG�Ͻ5�Ͻj�ϽP   P   ��Ͻ۱Ͻ��Ͻw�Ͻ��Ͻ�ϽW�Ͻ�Ͻw�ϽǱϽ�Ͻ	�ϽC�Ͻ��Ͻ.�Ͻ&�Ͻe�Ͻn�Ͻj�ϽӱϽP   P   ӱϽ̱Ͻ��Ͻ��Ͻp�Ͻs�Ͻ�Ͻ.�ϽױϽѱϽ�ϽڱϽ�Ͻ�ϽA�Ͻ'�Ͻv�Ͻ��Ͻ�Ͻ��ϽP   P   j�ϽαϽw�Ͻ�Ͻ̱Ͻ/�ϽN�Ͻ#�Ͻ
�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ߱Ͻ�Ͻ9�Ͻ3�Ͻt�Ͻ�ϽP   P   n�Ͻt�Ͻn�Ͻo�Ͻy�Ͻ�Ͻ3�Ͻ��Ͻ=�Ͻf�Ͻ�Ͻw�Ͻ��Ͻ�Ͻ|�ϽU�Ͻ��Ͻ:�Ͻ3�Ͻ��ϽP   P   e�ϽO�Ͻ�Ͻ,�Ͻ��Ͻ��Ͻa�Ͻ��ϽұϽ��Ͻ0�Ͻ��Ͻ1�Ͻo�Ͻ4�Ͻ��Ͻ��Ͻ��Ͻ9�Ͻv�ϽP   P   &�Ͻ��Ͻ2�Ͻ\�ϽO�Ͻ�Ͻ'�Ͻ�Ͻ>�Ͻ��Ͻ��Ͻ+�Ͻ�Ͻ��ϽM�Ͻ��Ͻ��ϽU�Ͻ�Ͻ'�ϽP   P   .�Ͻ˱Ͻ�Ͻ��Ͻ.�ϽڱϽD�Ͻ>�Ͻ�Ͻ��Ͻ�ϽN�Ͻ*�Ͻ��Ͻ��ϽM�Ͻ4�Ͻ|�Ͻ߱ϽA�ϽP   P   ��ϽN�Ͻ�Ͻ��ϽJ�Ͻ$�Ͻ:�ϽǲϽ��Ͻ�Ͻ+�Ͻm�Ͻ��Ͻw�Ͻ��Ͻ��Ͻo�Ͻ�Ͻ�Ͻ�ϽP   P   C�ϽE�Ͻ��ϽT�ϽO�Ͻ��Ͻ�Ͻ9�ϽM�Ͻ��Ͻ��Ͻ��Ͻ?�Ͻ��Ͻ*�Ͻ�Ͻ1�Ͻ��Ͻ��Ͻ�ϽP   P   	�Ͻ4�Ͻ �Ͻ��Ͻm�Ͻw�Ͻ[�ϽR�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻm�ϽN�Ͻ+�Ͻ��Ͻw�Ͻ��ϽڱϽP   P   �Ͻm�Ͻ�Ͻ�ϽV�ϽH�Ͻs�Ͻ�ϽX�Ͻv�Ͻ
�Ͻ��Ͻ��Ͻ+�Ͻ�Ͻ��Ͻ0�Ͻ�Ͻ��Ͻ�ϽP   P   ǱϽ|�Ͻ?�Ͻu�Ͻy�Ͻj�ϽN�Ͻ��Ͻc�ϽY�Ͻv�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻf�Ͻ�ϽѱϽP   P   w�Ͻ@�Ͻ|�Ͻ\�Ͻy�Ͻm�Ͻ��Ͻg�Ͻx�Ͻc�ϽX�Ͻ�ϽM�Ͻ��Ͻ�Ͻ>�ϽұϽ=�Ͻ
�ϽױϽP   P   �Ͻ�Ͻ	�Ͻ�Ͻ��Ͻ{�Ͻ��Ͻ�Ͻg�Ͻ��Ͻ�ϽR�Ͻ9�ϽǲϽ>�Ͻ�Ͻ��Ͻ��Ͻ#�Ͻ.�ϽP   P   W�Ͻ)�ϽW�Ͻ~�Ͻf�ϽG�Ͻ"�Ͻ��Ͻ��ϽN�Ͻs�Ͻ[�Ͻ�Ͻ:�ϽD�Ͻ'�Ͻa�Ͻ3�ϽN�Ͻ�ϽP   P   �ϽرϽ�Ͻ%�ϽO�Ͻr�ϽG�Ͻ{�Ͻm�Ͻj�ϽH�Ͻw�Ͻ��Ͻ$�ϽڱϽ�Ͻ��Ͻ�Ͻ/�Ͻs�ϽP   P   ��ϽO�ϽV�Ͻg�Ͻ��ϽO�Ͻf�Ͻ��Ͻy�Ͻy�ϽV�Ͻm�ϽO�ϽJ�Ͻ.�ϽO�Ͻ��Ͻy�Ͻ̱Ͻp�ϽP   P   w�Ͻ'�ϽL�Ͻ��Ͻg�Ͻ%�Ͻ~�Ͻ�Ͻ\�Ͻu�Ͻ�Ͻ��ϽT�Ͻ��Ͻ��Ͻ\�Ͻ,�Ͻo�Ͻ�Ͻ��ϽP   P   ��Ͻo�Ͻ�ϽL�ϽV�Ͻ�ϽW�Ͻ	�Ͻ|�Ͻ?�Ͻ�Ͻ �Ͻ��Ͻ�Ͻ�Ͻ2�Ͻ�Ͻn�Ͻw�Ͻ��ϽP   P   ۱ϽǱϽo�Ͻ'�ϽO�ϽرϽ)�Ͻ�Ͻ@�Ͻ|�Ͻm�Ͻ4�ϽE�ϽN�Ͻ˱Ͻ��ϽO�Ͻu�ϽαϽ̱ϽP   P   4�Ͻ��Ͻ5�Ͻ�ϽC�Ͻ1�ϽG�Ͻ��Ͻ��Ͻt�Ͻ��Ͻ��ϽB�ϽճϽ(�ϽN�Ͻ׳Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ|�Ͻ_�Ͻ�Ͻi�Ͻ˳Ͻb�ϽF�Ͻ�Ͻ��Ͻ��Ͻ��Ͻy�Ͻs�ϽJ�Ͻx�Ͻ�Ͻ��Ͻ1�ϽC�ϽP   P   �Ͻ��Ͻ �Ͻ2�Ͻ�Ͻ&�Ͻ��Ͻ��Ͻn�Ͻj�Ͻ6�Ͻ!�ϽH�Ͻ<�Ͻ?�Ͻ��ϽP�Ͻ�Ͻ��Ͻ1�ϽP   P   ��Ͻ�Ͻ'�Ͻ�Ͻy�Ͻ۳Ͻ,�Ͻ��Ͻ`�Ͻ$�Ͻ��Ͻ�ϽӳϽ��Ͻ&�Ͻ|�Ͻ��ϽE�Ͻ�Ͻ��ϽP   P   ׳Ͻ=�Ͻk�ϽE�Ͻ�Ͻ�Ͻh�Ͻ��ϽN�Ͻ=�Ͻ\�Ͻ��Ͻ˳ϽT�Ͻc�Ͻ0�Ͻ�Ͻ��ϽP�Ͻ�ϽP   P   N�Ͻ�Ͻ�Ͻ)�Ͻ�Ͻ(�Ͻn�Ͻ��ϽZ�Ͻ"�Ͻ��ϽE�ϽW�Ͻ��Ͻl�Ͻ�Ͻ0�Ͻ|�Ͻ��Ͻx�ϽP   P   (�Ͻs�Ͻ�Ͻ~�Ͻ�Ͻ��Ͻ�Ͻ`�Ͻ\�ϽW�ϽG�Ͻs�Ͻ��ϽʹϽL�Ͻl�Ͻc�Ͻ&�Ͻ?�ϽJ�ϽP   P   ճϽd�Ͻ�Ͻh�Ͻ@�Ͻl�ϽK�ϽݳϽ_�Ͻ�Ͻ�ϽT�Ͻ��Ͻ��ϽʹϽ��ϽT�Ͻ��Ͻ<�Ͻs�ϽP   P   B�ϽD�Ͻw�Ͻ��Ͻ�Ͻ.�Ͻd�Ͻl�Ͻ/�Ͻ��Ͻ'�Ͻ׳Ͻ�Ͻ��Ͻ��ϽW�Ͻ˳ϽӳϽH�Ͻy�ϽP   P   ��Ͻg�Ͻl�ϽS�Ͻ2�Ͻ'�Ͻ�Ͻ��ϽT�Ͻ��Ͻ��Ͻ�Ͻ׳ϽT�Ͻs�ϽE�Ͻ��Ͻ�Ͻ!�Ͻ��ϽP   P   ��Ͻ�Ͻ��ϽͳϽ��ϽY�Ͻ �Ͻ�ϽӳϽD�Ͻk�Ͻ��Ͻ'�Ͻ�ϽG�Ͻ��Ͻ\�Ͻ��Ͻ6�Ͻ��ϽP   P   t�ϽD�Ͻ!�Ͻ^�Ͻ�Ͻ��ϽZ�Ͻ�Ͻ:�Ͻ?�ϽD�Ͻ��Ͻ��Ͻ�ϽW�Ͻ"�Ͻ=�Ͻ$�Ͻj�Ͻ��ϽP   P   ��ϽL�Ͻ�Ͻ�Ͻ8�Ͻ�Ͻw�Ͻ(�Ͻ.�Ͻ:�ϽӳϽT�Ͻ/�Ͻ_�Ͻ\�ϽZ�ϽN�Ͻ`�Ͻn�Ͻ�ϽP   P   ��Ͻ-�ϽP�Ͻ��Ͻ�ϽS�ϽдϽ!�Ͻ(�Ͻ�Ͻ�Ͻ��Ͻl�ϽݳϽ`�Ͻ��Ͻ��Ͻ��Ͻ��ϽF�ϽP   P   G�Ͻ�Ͻ�Ͻ�Ͻ$�Ͻ0�Ͻ��ϽдϽw�ϽZ�Ͻ �Ͻ�Ͻd�ϽK�Ͻ�Ͻn�Ͻh�Ͻ,�Ͻ��Ͻb�ϽP   P   1�Ͻ��Ͻg�Ͻ�Ͻ�Ͻ��Ͻ0�ϽS�Ͻ�Ͻ��ϽY�Ͻ'�Ͻ.�Ͻl�Ͻ��Ͻ(�Ͻ�Ͻ۳Ͻ&�Ͻ˳ϽP   P   C�Ͻ��ϽL�Ͻ1�Ͻ��Ͻ�Ͻ$�Ͻ�Ͻ8�Ͻ�Ͻ��Ͻ2�Ͻ�Ͻ@�Ͻ�Ͻ�Ͻ�Ͻy�Ͻ�Ͻi�ϽP   P   �Ͻ��Ͻ'�Ͻh�Ͻ1�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ^�ϽͳϽS�Ͻ��Ͻh�Ͻ~�Ͻ)�ϽE�Ͻ�Ͻ2�Ͻ�ϽP   P   5�Ͻ�Ͻ��Ͻ'�ϽL�Ͻg�Ͻ�ϽP�Ͻ�Ͻ!�Ͻ��Ͻl�Ͻw�Ͻ�Ͻ�Ͻ�Ͻk�Ͻ'�Ͻ �Ͻ_�ϽP   P   ��Ͻ,�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ-�ϽL�ϽD�Ͻ�Ͻg�ϽD�Ͻd�Ͻs�Ͻ�Ͻ=�Ͻ�Ͻ��Ͻ|�ϽP   P   �Ͻ�ϽP�Ͻr�Ͻw�Ͻ��ϽV�Ͻg�Ͻ*�Ͻ��Ͻ��Ͻ�Ͻ�ϽM�Ͻ9�Ͻ��ϽC�Ͻz�Ͻ.�Ͻ�ϽP   P   �Ͻ�Ͻ�ϽR�Ͻ�Ͻ,�Ͻ%�Ͻ:�Ͻ\�Ͻ�Ͻ�Ͻ��Ͻ
�Ͻ��Ͻ4�Ͻ+�ϽP�Ͻ�Ͻp�Ͻ�ϽP   P   .�Ͻx�Ͻ@�Ͻi�ϽH�Ͻs�Ͻ0�Ͻ��ϽO�Ͻ��Ͻ"�Ͻ�Ͻ#�Ͻ��Ͻ<�Ͻ��Ͻ��Ͻl�Ͻ+�Ͻp�ϽP   P   z�Ͻ4�Ͻ)�ϽW�Ͻ��Ͻ]�ϽG�Ͻ�Ͻ�Ͻ�Ͻ~�Ͻ�ϽʶϽ��Ͻ(�Ͻ�Ͻ$�ϽP�Ͻl�Ͻ�ϽP   P   C�Ͻ��Ͻ<�Ͻ��ϽG�ϽZ�Ͻ�Ͻ/�Ͻ��Ͻ�Ͻt�Ͻ8�Ͻn�Ͻ�ϽI�Ͻ�Ͻs�Ͻ$�Ͻ��ϽP�ϽP   P   ��Ͻq�ϽN�ϽB�Ͻ_�Ͻ��Ͻ/�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�Ͻ�ϽB�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��Ͻ+�ϽP   P   9�Ͻq�Ͻ0�Ͻ��Ͻ1�Ͻ��Ͻ8�Ͻ>�ϽD�Ͻ/�Ͻd�Ͻ��Ͻ��Ͻ�Ͻv�Ͻ��ϽI�Ͻ(�Ͻ<�Ͻ4�ϽP   P   M�Ͻ?�ϽI�Ͻ�Ͻ�Ͻ:�Ͻ$�ϽH�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�ϽB�Ͻ�Ͻ��Ͻ��Ͻ��ϽP   P   �Ͻ7�Ͻ�ϽJ�Ͻ��Ͻd�Ͻ'�ϽQ�Ͻ��Ͻ�Ͻ1�ϽֶϽ��Ͻ�Ͻ��Ͻ�Ͻn�ϽʶϽ#�Ͻ
�ϽP   P   �Ͻm�ϽZ�Ͻt�Ͻ��Ͻ��Ͻk�ϽL�ϽN�Ͻ�Ͻ��Ͻ�ϽֶϽ��Ͻ��Ͻ�Ͻ8�Ͻ�Ͻ�Ͻ��ϽP   P   ��Ͻ0�Ͻ}�ϽL�Ͻ��Ͻ�Ͻ��Ͻa�Ͻ��Ͻ6�ϽڵϽ��Ͻ1�Ͻ��Ͻd�Ͻ�Ͻt�Ͻ~�Ͻ"�Ͻ�ϽP   P   ��Ͻ;�Ͻ��Ͻ��Ͻ��Ͻj�ϽU�Ͻ��Ͻ�Ͻ��Ͻ6�Ͻ�Ͻ�Ͻ��Ͻ/�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�ϽP   P   *�ϽL�Ͻ��Ͻr�Ͻu�Ͻ5�Ͻ��Ͻ8�Ͻ��Ͻ�Ͻ��ϽN�Ͻ��Ͻ��ϽD�Ͻ�Ͻ��Ͻ�ϽO�Ͻ\�ϽP   P   g�Ͻ<�Ͻ?�Ͻb�Ͻ��Ͻd�ϽߵϽ��Ͻ8�Ͻ��Ͻa�ϽL�ϽQ�ϽH�Ͻ>�Ͻ��Ͻ/�Ͻ�Ͻ��Ͻ:�ϽP   P   V�Ͻ�ϽM�ϽT�Ͻ��ϽK�Ͻ�ϽߵϽ��ϽU�Ͻ��Ͻk�Ͻ'�Ͻ$�Ͻ8�Ͻ/�Ͻ�ϽG�Ͻ0�Ͻ%�ϽP   P   ��Ͻ��ϽL�ϽK�Ͻz�Ͻ0�ϽK�Ͻd�Ͻ5�Ͻj�Ͻ�Ͻ��Ͻd�Ͻ:�Ͻ��Ͻ��ϽZ�Ͻ]�Ͻs�Ͻ,�ϽP   P   w�Ͻk�Ͻ:�Ͻ�ϽŶϽz�Ͻ��Ͻ��Ͻu�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ1�Ͻ_�ϽG�Ͻ��ϽH�Ͻ�ϽP   P   r�Ͻg�Ͻ8�Ͻ �Ͻ�ϽK�ϽT�Ͻb�Ͻr�Ͻ��ϽL�Ͻt�ϽJ�Ͻ�Ͻ��ϽB�Ͻ��ϽW�Ͻi�ϽR�ϽP   P   P�Ͻ5�Ͻr�Ͻ8�Ͻ:�ϽL�ϽM�Ͻ?�Ͻ��Ͻ��Ͻ}�ϽZ�Ͻ�ϽI�Ͻ0�ϽN�Ͻ<�Ͻ)�Ͻ@�Ͻ�ϽP   P   �ϽY�Ͻ5�Ͻg�Ͻk�Ͻ��Ͻ�Ͻ<�ϽL�Ͻ;�Ͻ0�Ͻm�Ͻ7�Ͻ?�Ͻq�Ͻq�Ͻ��Ͻ4�Ͻx�Ͻ�ϽP   P   �ϽD�ϽM�ϽX�Ͻ7�Ͻ�Ͻ�Ͻ��Ͻ3�Ͻ��Ͻj�Ͻh�ϽW�Ͻ��Ͻ*�Ͻ�ϽX�Ͻe�ϽK�ϽD�ϽP   P   D�Ͻ]�Ͻg�Ͻ��Ͻ+�Ͻ��Ͻq�Ͻj�Ͻ�ϽF�ϽԸϽ�Ͻp�ϽŷϽe�ϽZ�Ͻ��Ͻ�Ͻd�Ͻ��ϽP   P   K�Ͻ(�Ͻp�Ͻa�Ͻ��ϽK�Ͻ��Ͻ��ϽO�ϽշϽ"�Ͻu�Ͻ�ϽƷϽ_�Ͻ��Ͻ��Ͻh�ϽַϽd�ϽP   P   e�ϽT�Ͻ&�Ͻw�Ͻ!�Ͻz�Ͻ%�Ͻ:�Ͻ�ϽX�Ͻ!�Ͻ�Ͻ�Ͻ?�Ͻ{�Ͻ��Ͻ3�Ͻ�Ͻh�Ͻ�ϽP   P   X�Ͻ��Ͻ�Ͻ�ϽY�Ͻ��Ͻy�Ͻ�Ͻ��Ͻ2�Ͻ�Ͻ�Ͻ�Ͻ�Ͻ�ϽB�Ͻ��Ͻ3�Ͻ��Ͻ��ϽP   P   �Ͻ�Ͻ[�ϽZ�Ͻ�Ͻ��ϽY�ϽʸϽ۸ϽA�Ͻ0�Ͻi�Ͻ��Ͻ��Ͻ��ϽM�ϽB�Ͻ��Ͻ��ϽZ�ϽP   P   *�ϽķϽ��Ͻ��Ͻ��Ͻ÷Ͻ<�ϽQ�ϽR�ϽC�Ͻ+�Ͻo�Ͻ�ϽO�ϽθϽ��Ͻ�Ͻ{�Ͻ_�Ͻe�ϽP   P   ��ϽN�ϽJ�Ͻq�Ͻ��Ͻ8�Ͻ?�ϽøϽ޷Ͻ�Ͻ�Ͻ�Ͻ��ϽB�ϽO�Ͻ��Ͻ�Ͻ?�ϽƷϽŷϽP   P   W�Ͻe�Ͻ8�Ͻb�Ͻ5�Ͻ9�ϽX�Ͻk�Ͻo�Ͻ.�Ͻ=�Ͻ��Ͻ0�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�Ͻ�Ͻp�ϽP   P   h�Ͻ3�Ͻ#�Ͻ%�Ͻ��Ͻ�Ͻ:�Ͻ�Ͻ5�Ͻ��Ͻ��Ͻp�Ͻ��Ͻ�Ͻo�Ͻi�Ͻ�Ͻ�Ͻu�Ͻ�ϽP   P   j�Ͻ��Ͻ*�ϽX�Ͻ@�Ͻ�ϽG�ϽD�Ͻt�ϽP�Ͻ��Ͻ��Ͻ=�Ͻ�Ͻ+�Ͻ0�Ͻ�Ͻ!�Ͻ"�ϽԸϽP   P   ��ϽV�ϽڷϽϷϽ/�Ͻ�Ͻ9�Ͻ�ϽѷϽƷϽP�Ͻ��Ͻ.�Ͻ�ϽC�ϽA�Ͻ2�ϽX�ϽշϽF�ϽP   P   3�ϽR�Ͻ1�Ͻ�Ͻ��Ͻz�Ͻ��Ͻ~�Ͻ*�ϽѷϽt�Ͻ5�Ͻo�Ͻ޷ϽR�Ͻ۸Ͻ��Ͻ�ϽO�Ͻ�ϽP   P   ��Ͻq�Ͻ1�ϽF�Ͻ �Ͻr�Ͻ��Ͻl�Ͻ~�Ͻ�ϽD�Ͻ�Ͻk�ϽøϽQ�ϽʸϽ�Ͻ:�Ͻ��Ͻj�ϽP   P   �Ͻc�Ͻ�ϽG�Ͻ.�ϽM�Ͻu�Ͻ��Ͻ��Ͻ9�ϽG�Ͻ:�ϽX�Ͻ?�Ͻ<�ϽY�Ͻy�Ͻ%�Ͻ��Ͻq�ϽP   P   �ϽŷϽN�Ͻc�Ͻ�Ͻ�ϽM�Ͻr�Ͻz�Ͻ�Ͻ�Ͻ�Ͻ9�Ͻ8�Ͻ÷Ͻ��Ͻ��Ͻz�ϽK�Ͻ��ϽP   P   7�Ͻ�Ͻ_�Ͻ��Ͻ�Ͻ�Ͻ.�Ͻ �Ͻ��Ͻ/�Ͻ@�Ͻ��Ͻ5�Ͻ��Ͻ��Ͻ�ϽY�Ͻ!�Ͻ��Ͻ+�ϽP   P   X�Ͻ&�Ͻ\�ϽָϽ��Ͻc�ϽG�ϽF�Ͻ�ϽϷϽX�Ͻ%�Ͻb�Ͻq�Ͻ��ϽZ�Ͻ�Ͻw�Ͻa�Ͻ��ϽP   P   M�Ͻ7�Ͻ߷Ͻ\�Ͻ_�ϽN�Ͻ�Ͻ1�Ͻ1�ϽڷϽ*�Ͻ#�Ͻ8�ϽJ�Ͻ��Ͻ[�Ͻ�Ͻ&�Ͻp�Ͻg�ϽP   P   D�Ͻ@�Ͻ7�Ͻ&�Ͻ�ϽŷϽc�Ͻq�ϽR�ϽV�Ͻ��Ͻ3�Ͻe�ϽN�ϽķϽ�Ͻ��ϽT�Ͻ(�Ͻ]�ϽP   P   	�Ͻ7�Ͻ��Ͻ�Ͻ�Ͻ��ϽR�Ͻ˹Ͻ�Ͻ9�Ͻ��Ͻ�ϽV�Ͻ�Ͻ��Ͻ��Ͻy�Ͻ��Ͻ�Ͻ1�ϽP   P   1�ϽN�Ͻ9�Ͻ1�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��ϽֹϽ޺ϽN�Ͻ�Ͻ��ϽʹϽz�Ͻ�Ͻk�ϽP   P   �Ͻ=�Ͻ�Ͻ�Ͻ��Ͻ�ϽҹϽ1�Ͻ�Ͻ��ϽZ�Ͻ<�Ͻ4�Ͻ�ϽL�ϽB�Ͻ�Ͻ�Ͻ�Ͻ�ϽP   P   ��Ͻ��Ͻg�Ͻ��Ͻ��Ͻ>�Ͻ�Ͻr�Ͻ�ϽP�Ͻ��Ͻ4�Ͻ5�Ͻ��ϽW�Ͻ��ϽN�ϽE�Ͻ�Ͻz�ϽP   P   y�Ͻ'�ϽǺϽ=�Ͻ]�Ͻ��Ͻ��Ͻ(�Ͻ��Ͻ@�Ͻs�Ͻ��Ͻo�ϽѺϽW�ϽH�Ͻ�ϽN�Ͻ�ϽʹϽP   P   ��Ͻ��ϽG�Ͻ=�Ͻ��Ͻ��Ͻ�Ͻ^�Ͻ��Ͻg�Ͻ�Ͻ-�Ͻ�ϽչϽ�Ͻ�ϽH�Ͻ��ϽB�Ͻ��ϽP   P   ��ϽͺϽG�Ͻ��ϽL�ϽʺϽ��Ͻ��Ͻ"�Ͻ#�Ͻ��Ͻ�Ͻ	�Ͻ�Ͻ=�Ͻ�ϽW�ϽW�ϽL�Ͻ�ϽP   P   �Ͻ+�ϽE�Ͻ�Ͻ�ϽG�Ͻ3�ϽԹϽa�Ͻ��Ͻw�ϽҺϽ�Ͻ�Ͻ�ϽչϽѺϽ��Ͻ�ϽN�ϽP   P   V�Ͻ"�Ͻ��ϽX�ϽK�Ͻ7�Ͻ��Ͻ�ϽZ�Ͻ��Ͻ[�Ͻ8�ϽW�Ͻ�Ͻ	�Ͻ�Ͻo�Ͻ5�Ͻ4�Ͻ޺ϽP   P   �Ͻ�Ͻz�Ͻ,�Ͻ}�Ͻy�Ͻg�ϽG�Ͻ �Ͻ�ϽùϽ?�Ͻ8�ϽҺϽ�Ͻ-�Ͻ��Ͻ4�Ͻ<�ϽֹϽP   P   ��Ͻ��ϽW�Ͻu�ϽU�Ͻ�ϽG�ϽX�Ͻ��ϽS�Ͻ�ϽùϽ[�Ͻw�Ͻ��Ͻ�Ͻs�Ͻ��ϽZ�Ͻ��ϽP   P   9�ϽF�Ͻ@�Ͻ˺Ͻ=�Ͻ*�ϽT�Ͻ�ϽںϽ.�ϽS�Ͻ�Ͻ��Ͻ��Ͻ#�Ͻg�Ͻ@�ϽP�Ͻ��Ͻ��ϽP   P   �Ͻ)�ϽL�Ͻ�Ͻ��Ͻ+�ϽN�Ͻ�Ͻ��ϽںϽ��Ͻ �ϽZ�Ͻa�Ͻ"�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��ϽP   P   ˹Ͻ7�Ͻ��Ͻ9�Ͻ(�Ͻ�Ͻ8�Ͻ�Ͻ�Ͻ�ϽX�ϽG�Ͻ�ϽԹϽ��Ͻ^�Ͻ(�Ͻr�Ͻ1�Ͻ�ϽP   P   R�Ͻx�Ͻ>�Ͻ]�Ͻ7�Ͻu�Ͻ�Ͻ8�ϽN�ϽT�ϽG�Ͻg�Ͻ��Ͻ3�Ͻ��Ͻ�Ͻ��Ͻ�ϽҹϽ�ϽP   P   ��ϽܺϽ\�Ͻ}�Ͻ��ϽܺϽu�Ͻ�Ͻ+�Ͻ*�Ͻ�Ͻy�Ͻ7�ϽG�ϽʺϽ��Ͻ��Ͻ>�Ͻ�Ͻ�ϽP   P   �Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ7�Ͻ(�Ͻ��Ͻ=�ϽU�Ͻ}�ϽK�Ͻ�ϽL�Ͻ��Ͻ]�Ͻ��Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻ6�Ͻ¹Ͻ�Ͻ}�Ͻ]�Ͻ9�Ͻ�Ͻ˺Ͻu�Ͻ,�ϽX�Ͻ�Ͻ��Ͻ=�Ͻ=�Ͻ��Ͻ�Ͻ1�ϽP   P   ��Ͻ��Ͻp�Ͻ6�Ͻ��Ͻ\�Ͻ>�Ͻ��ϽL�Ͻ@�ϽW�Ͻz�Ͻ��ϽE�ϽG�ϽG�ϽǺϽg�Ͻ�Ͻ9�ϽP   P   7�Ͻb�Ͻ��Ͻ��Ͻ��ϽܺϽx�Ͻ7�Ͻ)�ϽF�Ͻ��Ͻ�Ͻ"�Ͻ+�ϽͺϽ��Ͻ'�Ͻ��Ͻ=�ϽN�ϽP   P   �Ͻ]�Ͻ��Ͻy�Ͻ�Ͻ+�Ͻ(�ϽE�ϽJ�Ͻt�Ͻ��Ͻ<�Ͻu�ϽQ�Ͻj�Ͻ�Ͻh�Ͻ��Ͻ��ϽT�ϽP   P   T�ϽP�Ͻ~�Ͻ�Ͻu�Ͻ��Ͻ��Ͻ��Ͻ��ϽλϽD�Ͻ��ϽлϽf�Ͻf�Ͻn�Ͻe�ϽC�Ͻ$�Ͻo�ϽP   P   ��ϽM�Ͻ��ϽA�Ͻ �Ͻ%�ϽL�Ͻ=�ϽM�Ͻ�Ͻ7�ϽݼϽ8�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ3�ϽT�Ͻ$�ϽP   P   ��Ͻ�Ͻ"�Ͻ~�Ͻb�Ͻ-�Ͻ��Ͻ��Ͻ9�ϽM�Ͻ�Ͻ@�Ͻ)�Ͻ�Ͻ�Ͻ+�Ͻm�Ͻ[�Ͻ3�ϽC�ϽP   P   h�Ͻ)�Ͻ�ϽB�Ͻ;�Ͻ��Ͻi�Ͻi�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ9�Ͻ'�Ͻ��ϽμϽm�Ͻ��Ͻe�ϽP   P   �Ͻ�Ͻn�ϽF�Ͻ�Ͻ�Ͻ��Ͻ5�ϽK�Ͻ��Ͻz�Ͻ~�Ͻ<�Ͻ�Ͻ8�Ͻ��Ͻ��Ͻ+�Ͻ�Ͻn�ϽP   P   j�Ͻ�ϽV�Ͻ��Ͻ:�Ͻ�Ͻ@�Ͻ��ϽJ�Ͻ�Ͻ�ϽR�Ͻ?�Ͻ��Ͻ��Ͻ8�Ͻ'�Ͻ�Ͻ��Ͻf�ϽP   P   Q�Ͻ�Ͻ�Ͻ��ϽռϽ��Ͻ&�ϽZ�Ͻt�Ͻ@�Ͻ�ϽM�Ͻ:�Ͻ�Ͻ��Ͻ�Ͻ9�Ͻ�Ͻ�Ͻf�ϽP   P   u�Ͻo�ϽC�Ͻ0�Ͻ��Ͻ�Ͻ,�Ͻ�Ͻ^�ϽܻϽ�ϽN�Ͻ?�Ͻ:�Ͻ?�Ͻ<�Ͻ��Ͻ)�Ͻ8�ϽлϽP   P   <�Ͻ`�Ͻ@�Ͻ �Ͻ�Ͻ�ϽH�Ͻ,�Ͻt�ϽG�Ͻ~�ϽټϽN�ϽM�ϽR�Ͻ~�Ͻ�Ͻ@�ϽݼϽ��ϽP   P   ��Ͻo�Ͻ�Ͻ+�Ͻ=�ϽλϽ-�Ͻ)�Ͻ�Ͻl�Ͻ߼Ͻ~�Ͻ�Ͻ�Ͻ�Ͻz�Ͻ��Ͻ�Ͻ7�ϽD�ϽP   P   t�Ͻ[�Ͻ�Ͻ�Ͻg�Ͻ7�ϽO�Ͻp�Ͻ��Ͻ��Ͻl�ϽG�ϽܻϽ@�Ͻ�Ͻ��Ͻ��ϽM�Ͻ�ϽλϽP   P   J�ϽB�Ͻ)�Ͻ �Ͻ �Ͻv�ϽD�Ͻ��Ͻ��Ͻ��Ͻ�Ͻt�Ͻ^�Ͻt�ϽJ�ϽK�Ͻ��Ͻ9�ϽM�Ͻ��ϽP   P   E�Ͻ��Ͻh�Ͻ�Ͻj�Ͻs�Ͻb�Ͻ[�Ͻ��Ͻp�Ͻ)�Ͻ,�Ͻ�ϽZ�Ͻ��Ͻ5�Ͻi�Ͻ��Ͻ=�Ͻ��ϽP   P   (�Ͻ/�Ͻ��Ͻ�ϽW�ϽI�Ͻ?�Ͻb�ϽD�ϽO�Ͻ-�ϽH�Ͻ,�Ͻ&�Ͻ@�Ͻ��Ͻi�Ͻ��ϽL�Ͻ��ϽP   P   +�Ͻ�Ͻ�ϽV�Ͻ�Ͻ��ϽI�Ͻs�Ͻv�Ͻ7�ϽλϽ�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ-�Ͻ%�Ͻ��ϽP   P   �Ͻ�Ͻ"�Ͻ��ϽN�Ͻ�ϽW�Ͻj�Ͻ �Ͻg�Ͻ=�Ͻ�Ͻ��ϽռϽ:�Ͻ�Ͻ;�Ͻb�Ͻ �Ͻu�ϽP   P   y�Ͻh�Ͻc�ϽʼϽ��ϽV�Ͻ�Ͻ�Ͻ �Ͻ�Ͻ+�Ͻ �Ͻ0�Ͻ��Ͻ��ϽF�ϽB�Ͻ~�ϽA�Ͻ�ϽP   P   ��Ͻ"�Ͻ̻Ͻc�Ͻ"�Ͻ�Ͻ��Ͻh�Ͻ)�Ͻ�Ͻ�Ͻ@�ϽC�Ͻ�ϽV�Ͻn�Ͻ�Ͻ"�Ͻ��Ͻ~�ϽP   P   ]�Ͻ1�Ͻ"�Ͻh�Ͻ�Ͻ�Ͻ/�Ͻ��ϽB�Ͻ[�Ͻo�Ͻ`�Ͻo�Ͻ�Ͻ�Ͻ�Ͻ)�Ͻ�ϽM�ϽP�ϽP   P   �Ͻ@�ϽN�ϽX�Ͻ@�Ͻ-�Ͻ&�Ͻ]�Ͻ]�Ͻq�Ͻ)�Ͻh�ϽY�ϽW�Ͻ9�Ͻ4�Ͻ;�ϽY�ϽA�ϽF�ϽP   P   F�Ͻ)�Ͻ��Ͻ;�Ͻ��Ͻo�Ͻ'�Ͻ&�Ͻ�Ͻe�Ͻ&�ϽK�Ͻ)�Ͻ
�Ͻ$�Ͻ&�Ͻn�ϽҽϽg�Ͻ�ϽP   P   A�Ͻ'�Ͻ!�Ͻy�Ͻ4�Ͻm�Ͻ;�Ͻ8�ϽG�ϽG�Ͻ��Ͻ߽Ͻ��ϽQ�ϽV�Ͻ'�ϽY�ϽY�Ͻ;�Ͻg�ϽP   P   Y�Ͻ.�ϽX�Ͻ?�Ͻ�ϽH�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻj�Ͻ��Ͻ�ϽɽϽY�ϽҽϽP   P   ;�Ͻv�Ͻ-�Ͻ{�Ͻ�Ͻ��Ͻ+�Ͻ��Ͻ�Ͻ��Ͻ!�Ͻ�ϽU�Ͻ�ϽP�Ͻ��Ͻ�Ͻ�ϽY�Ͻn�ϽP   P   4�ϽP�Ͻd�ϽF�Ͻ��Ͻ!�Ͻ'�Ͻ3�Ͻ��Ͻ��Ͻ�Ͻ��Ͻt�Ͻ{�Ͻg�Ͻ"�Ͻ��Ͻ��Ͻ'�Ͻ&�ϽP   P   9�Ͻ^�Ͻ]�Ͻ�ϽQ�Ͻw�Ͻ�Ͻ?�Ͻ1�Ͻ��Ͻ!�Ͻz�Ͻ�Ͻ̽ϽC�Ͻg�ϽP�Ͻj�ϽV�Ͻ$�ϽP   P   W�Ͻ��Ͻ��ϽܽϽ��Ͻ��Ͻ��ϽZ�Ͻ�Ͻ_�Ͻ��Ͻ-�Ͻx�Ͻ�Ͻ̽Ͻ{�Ͻ�Ͻ��ϽQ�Ͻ
�ϽP   P   Y�Ͻ0�ϽJ�Ͻ0�Ͻ�ϽD�Ͻ/�Ͻ1�Ͻ.�Ͻl�ϽZ�Ͻ'�Ͻ�Ͻx�Ͻ�Ͻt�ϽU�Ͻ��Ͻ��Ͻ)�ϽP   P   h�Ͻ<�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ9�ϽL�ϽS�Ͻ[�Ͻ�Ͻ'�Ͻ-�Ͻz�Ͻ��Ͻ�Ͻ�Ͻ߽ϽK�ϽP   P   )�Ͻ��Ͻ��Ͻ[�Ͻx�Ͻ�Ͻp�ϽY�Ͻo�Ͻ��Ͻ�Ͻ[�ϽZ�Ͻ��Ͻ!�Ͻ�Ͻ!�Ͻ��Ͻ��Ͻ&�ϽP   P   q�Ͻ۽ϽʾϽb�Ͻb�Ͻ��Ͻb�Ͻu�Ͻs�ϽӾϽ��ϽS�Ͻl�Ͻ_�Ͻ��Ͻ��Ͻ��Ͻ��ϽG�Ͻe�ϽP   P   ]�Ͻ	�Ͻ��Ͻ=�Ͻ,�ϽO�Ͻ
�ϽG�Ͻ�Ͻs�Ͻo�ϽL�Ͻ.�Ͻ�Ͻ1�Ͻ��Ͻ�Ͻ��ϽG�Ͻ�ϽP   P   ]�Ͻ=�Ͻ8�ϽI�Ͻh�ϽA�ϽM�Ͻ|�ϽG�Ͻu�ϽY�Ͻ9�Ͻ1�ϽZ�Ͻ?�Ͻ3�Ͻ��Ͻ�Ͻ8�Ͻ&�ϽP   P   &�Ͻ��ϽT�Ͻd�Ͻ��ϽF�ϽM�ϽM�Ͻ
�Ͻb�Ͻp�Ͻ��Ͻ/�Ͻ��Ͻ�Ͻ'�Ͻ+�Ͻ�Ͻ;�Ͻ'�ϽP   P   -�Ͻr�Ͻ��Ͻ`�Ͻ�Ͻ%�ϽF�ϽA�ϽO�Ͻ��Ͻ�Ͻ��ϽD�Ͻ��Ͻw�Ͻ!�Ͻ��ϽH�Ͻm�Ͻo�ϽP   P   @�Ͻ[�Ͻe�ϽܽϽ��Ͻ�Ͻ��Ͻh�Ͻ,�Ͻb�Ͻx�Ͻ��Ͻ�Ͻ��ϽQ�Ͻ��Ͻ�Ͻ�Ͻ4�Ͻ��ϽP   P   X�Ͻb�ϽK�Ͻ�ϽܽϽ`�Ͻd�ϽI�Ͻ=�Ͻb�Ͻ[�Ͻ��Ͻ0�ϽܽϽ�ϽF�Ͻ{�Ͻ?�Ͻy�Ͻ;�ϽP   P   N�ϽJ�Ͻ@�ϽK�Ͻe�Ͻ��ϽT�Ͻ8�Ͻ��ϽʾϽ��Ͻ�ϽJ�Ͻ��Ͻ]�Ͻd�Ͻ-�ϽX�Ͻ!�Ͻ��ϽP   P   @�Ͻ�ϽJ�Ͻb�Ͻ[�Ͻr�Ͻ��Ͻ=�Ͻ	�Ͻ۽Ͻ��Ͻ<�Ͻ0�Ͻ��Ͻ^�ϽP�Ͻv�Ͻ.�Ͻ'�Ͻ)�ϽP   P   �Ͻ?�ϽA�Ͻ�Ͻ��Ͻ|�Ͻs�Ͻ:�ϽE�ϽG�Ͻ9�Ͻ��Ͻ!�Ͻ�Ͻ:�Ͻ��ϽM�Ͻ�Ͻ'�Ͻ8�ϽP   P   8�ϽT�ϽC�Ͻr�Ͻ7�Ͻ�Ͻ2�Ͻd�Ͻo�Ͻ��Ͻ�Ͻ�Ͻ}�Ͻ��Ͻ��Ͻ(�Ͻ�Ͻe�Ͻ}�ϽF�ϽP   P   '�Ͻ��Ͻ�Ͻ��Ͻ��Ͻg�Ͻd�ϽS�Ͻ4�Ͻ�Ͻ9�Ͻ�ϽE�Ͻ0�Ͻ�ϽT�Ͻ(�Ͻf�Ͻ�Ͻ}�ϽP   P   �Ͻp�Ͻx�Ͻ&�ϽA�ϽY�Ͻ��Ͻo�ϽC�Ͻ�Ͻ5�Ͻ��Ͻ��Ͻ)�Ͻ��Ͻa�Ͻ��Ͻ��Ͻf�Ͻe�ϽP   P   M�Ͻ4�Ͻq�Ͻ�ϽW�Ͻ/�Ͻ>�Ͻ��Ͻ}�Ͻ}�Ͻ��ϽA�ϽY�Ͻ5�Ͻ��Ͻ��Ͻ,�Ͻ��Ͻ(�Ͻ�ϽP   P   ��Ͻg�Ͻ!�Ͻ,�Ͻ^�Ͻ��Ͻ�Ͻ_�Ͻ�Ͻq�Ͻ��Ͻ�Ͻ7�Ͻ2�Ͻ�Ͻ��Ͻ��Ͻa�ϽT�Ͻ(�ϽP   P   :�ϽJ�Ͻ�ϽR�Ͻ�Ͻ8�ϽL�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��ϽK�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��ϽP   P   �Ͻ�Ͻ&�Ͻ��Ͻq�Ͻ,�Ͻ�Ͻ6�Ͻu�Ͻ
�Ͻ2�Ͻ+�Ͻ>�Ͻm�Ͻ��Ͻ2�Ͻ5�Ͻ)�Ͻ0�Ͻ��ϽP   P   !�Ͻ9�Ͻ�ϽP�Ͻt�Ͻ[�Ͻ�Ͻ�Ͻ<�Ͻ��Ͻ5�Ͻ��Ͻ`�Ͻ>�ϽK�Ͻ7�ϽY�Ͻ��ϽE�Ͻ}�ϽP   P   ��ϽV�ϽM�Ͻ:�ϽD�ϽT�Ͻ�Ͻ��ϽU�ϽQ�Ͻ�Ͻ'�Ͻ��Ͻ+�Ͻ��Ͻ�ϽA�Ͻ��Ͻ�Ͻ�ϽP   P   9�ϽR�ϽT�Ͻ�ϽտϽw�Ͻ�Ͻ�Ͻ%�Ͻp�Ͻ9�Ͻ�Ͻ5�Ͻ2�Ͻ��Ͻ��Ͻ��Ͻ5�Ͻ9�Ͻ�ϽP   P   G�Ͻ}�Ͻ2�Ͻ/�Ͻ��Ͻq�ϽM�Ͻ5�ϽA�Ͻ)�Ͻp�ϽQ�Ͻ��Ͻ
�Ͻ�Ͻq�Ͻ}�Ͻ�Ͻ�Ͻ��ϽP   P   E�ϽR�ϽJ�Ͻ&�Ͻ��Ͻ+�Ͻ�Ͻ#�Ͻ��ϽA�Ͻ%�ϽU�Ͻ<�Ͻu�Ͻ�Ͻ�Ͻ}�ϽC�Ͻ4�Ͻo�ϽP   P   :�Ͻ	�Ͻd�Ͻ�Ͻ,�Ͻ�Ͻ2�Ͻk�Ͻ#�Ͻ5�Ͻ�Ͻ��Ͻ�Ͻ6�Ͻ��Ͻ_�Ͻ��Ͻo�ϽS�Ͻd�ϽP   P   s�Ͻ��ϽP�Ͻ�Ͻ��ϽB�Ͻv�Ͻ2�Ͻ�ϽM�Ͻ�Ͻ�Ͻ�Ͻ�ϽL�Ͻ�Ͻ>�Ͻ��Ͻd�Ͻ2�ϽP   P   |�Ͻ:�Ͻ�Ͻ@�Ͻ/�Ͻ��ϽB�Ͻ�Ͻ+�Ͻq�Ͻw�ϽT�Ͻ[�Ͻ,�Ͻ8�Ͻ��Ͻ/�ϽY�Ͻg�Ͻ�ϽP   P   ��ϽT�ϽM�Ͻn�Ͻ��Ͻ/�Ͻ��Ͻ,�Ͻ��Ͻ��ϽտϽD�Ͻt�Ͻq�Ͻ�Ͻ^�ϽW�ϽA�Ͻ��Ͻ7�ϽP   P   �Ͻ�Ͻ�Ͻ:�Ͻn�Ͻ@�Ͻ�Ͻ�Ͻ&�Ͻ/�Ͻ�Ͻ:�ϽP�Ͻ��ϽR�Ͻ,�Ͻ�Ͻ&�Ͻ��Ͻr�ϽP   P   A�Ͻe�Ͻ��Ͻ�ϽM�Ͻ�ϽP�Ͻd�ϽJ�Ͻ2�ϽT�ϽM�Ͻ�Ͻ&�Ͻ�Ͻ!�Ͻq�Ͻx�Ͻ�ϽC�ϽP   P   ?�Ͻ��Ͻe�Ͻ�ϽT�Ͻ:�Ͻ��Ͻ	�ϽR�Ͻ}�ϽR�ϽV�Ͻ9�Ͻ�ϽJ�Ͻg�Ͻ4�Ͻp�Ͻ��ϽT�ϽP   P   ��Ͻe�Ͻ>�Ͻ{�Ͻ��Ͻ��Ͻf�ϽJ�Ͻ1�Ͻ��Ͻn�Ͻ)�Ͻ��Ͻ1�Ͻ*�Ͻ�Ͻ#�Ͻh�Ͻ8�Ͻr�ϽP   P   r�Ͻ��Ͻp�Ͻ�Ͻf�Ͻ�Ͻx�Ͻ�ϽR�Ͻ��Ͻ��Ͻ��Ͻ��Ͻl�Ͻb�Ͻv�ϽE�Ͻ��Ͻ��Ͻ��ϽP   P   8�Ͻ�Ͻ4�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ*�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ*�ϽN�Ͻ#�Ͻ�Ͻ��Ͻ��ϽP   P   h�Ͻ&�Ͻ�Ͻ��Ͻg�Ͻ
�Ͻ��Ͻ��Ͻ+�Ͻ%�Ͻ��Ͻ�ϽJ�Ͻ��Ͻk�Ͻ4�Ͻ.�Ͻ6�Ͻ�Ͻ��ϽP   P   #�Ͻ#�Ͻ-�Ͻ�ϽW�Ͻ*�Ͻc�Ͻ(�Ͻ@�Ͻ:�ϽM�Ͻg�Ͻ��Ͻ^�Ͻ�Ͻl�Ͻ��Ͻ.�Ͻ#�ϽE�ϽP   P   �Ͻ+�ϽQ�Ͻ��Ͻ�Ͻ+�ϽF�ϽA�Ͻ��ϽI�Ͻ��Ͻ�ϽI�Ͻ5�Ͻ��Ͻ��Ͻl�Ͻ4�ϽN�Ͻv�ϽP   P   *�Ͻ4�Ͻ7�Ͻ��ϽY�Ͻ�Ͻb�Ͻ'�Ͻ��Ͻt�Ͻ6�Ͻ\�Ͻ��ϽH�Ͻ��Ͻ��Ͻ�Ͻk�Ͻ*�Ͻb�ϽP   P   1�Ͻt�Ͻ�Ͻu�Ͻ7�ϽN�Ͻ]�ϽA�Ͻ:�Ͻ]�Ͻ��ϽQ�ϽJ�Ͻ��ϽH�Ͻ5�Ͻ^�Ͻ��Ͻ��Ͻl�ϽP   P   ��Ͻ��ϽS�ϽO�Ͻ�ϽB�Ͻl�Ͻ��ϽI�Ͻ��Ͻ.�Ͻ�Ͻ�ϽJ�Ͻ��ϽI�Ͻ��ϽJ�Ͻ��Ͻ��ϽP   P   )�Ͻ6�Ͻ-�Ͻe�Ͻ��Ͻ�Ͻ5�Ͻi�Ͻ,�Ͻ��Ͻ�Ͻ��Ͻ�ϽQ�Ͻ\�Ͻ�Ͻg�Ͻ�Ͻ��Ͻ��ϽP   P   n�Ͻs�Ͻ��Ͻ��Ͻr�ϽT�Ͻr�Ͻ��Ͻ	�Ͻu�Ͻ��Ͻ�Ͻ.�Ͻ��Ͻ6�Ͻ��ϽM�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ�Ͻ?�ϽN�Ͻ-�Ͻe�Ͻ �Ͻ�Ͻu�Ͻ��Ͻ��Ͻ]�Ͻt�ϽI�Ͻ:�Ͻ%�Ͻ��Ͻ��ϽP   P   1�Ͻg�Ͻ��Ͻ&�ϽS�Ͻ^�Ͻ��ϽB�Ͻ<�Ͻ �Ͻ	�Ͻ,�ϽI�Ͻ:�Ͻ��Ͻ��Ͻ@�Ͻ+�Ͻ��ϽR�ϽP   P   J�Ͻ��Ͻ7�Ͻ��Ͻ`�Ͻ#�ϽX�Ͻl�ϽB�Ͻe�Ͻ��Ͻi�Ͻ��ϽA�Ͻ'�ϽA�Ͻ(�Ͻ��Ͻ*�Ͻ�ϽP   P   f�Ͻ]�Ͻ��Ͻq�ϽM�Ͻ:�Ͻ��ϽX�Ͻ��Ͻ-�Ͻr�Ͻ5�Ͻl�Ͻ]�Ͻb�ϽF�Ͻc�Ͻ��Ͻ�Ͻx�ϽP   P   ��Ͻ�Ͻ/�Ͻ�Ͻ�Ͻo�Ͻ:�Ͻ#�Ͻ^�ϽN�ϽT�Ͻ�ϽB�ϽN�Ͻ�Ͻ+�Ͻ*�Ͻ
�Ͻ�Ͻ�ϽP   P   ��Ͻ�Ͻq�ϽU�ϽW�Ͻ�ϽM�Ͻ`�ϽS�Ͻ?�Ͻr�Ͻ��Ͻ�Ͻ7�ϽY�Ͻ�ϽW�Ͻg�Ͻ��Ͻf�ϽP   P   {�Ͻ��Ͻ`�Ͻo�ϽU�Ͻ�Ͻq�Ͻ��Ͻ&�Ͻ�Ͻ��Ͻe�ϽO�Ͻu�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�ϽP   P   >�Ͻ��Ͻy�Ͻ`�Ͻq�Ͻ/�Ͻ��Ͻ7�Ͻ��Ͻ��Ͻ��Ͻ-�ϽS�Ͻ�Ͻ7�ϽQ�Ͻ-�Ͻ�Ͻ4�Ͻp�ϽP   P   e�Ͻ6�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ]�Ͻ��Ͻg�Ͻ��Ͻs�Ͻ6�Ͻ��Ͻt�Ͻ4�Ͻ+�Ͻ#�Ͻ&�Ͻ�Ͻ��ϽP   P   ~�Ͻ�Ͻ6�ϽT�Ͻ�Ͻ1�Ͻ`�Ͻ4�Ͻ��ϽA�Ͻ��Ͻq�Ͻk�Ͻ+�Ͻ6�Ͻ,�Ͻ �ϽK�Ͻ7�Ͻ�ϽP   P   �Ͻ(�Ͻ�Ͻw�Ͻ�Ͻ>�ϽY�Ͻ��Ͻ�ϽM�Ͻ2�Ͻ�Ͻe�Ͻ�Ͻ �Ͻ^�Ͻ^�ϽK�Ͻf�Ͻ �ϽP   P   7�Ͻ�Ͻ:�Ͻ]�Ͻ��Ͻ��Ͻc�Ͻ�Ͻ5�Ͻ��ϽX�Ͻ��ϽQ�Ͻ��Ͻ��Ͻ4�Ͻ0�Ͻ��Ͻ��Ͻf�ϽP   P   K�Ͻ��Ͻ�ϽW�Ͻ:�Ͻ��Ͻ�ϽG�Ͻz�ϽB�Ͻ��Ͻ*�ϽU�Ͻ��Ͻb�Ͻ��ϽX�ϽJ�Ͻ��ϽK�ϽP   P    �Ͻ��ϽC�Ͻj�Ͻ�ϽG�Ͻt�Ͻf�Ͻq�Ͻ�ϽJ�Ͻ��ϽS�Ͻ��Ͻ-�Ͻ>�ϽK�ϽX�Ͻ0�Ͻ^�ϽP   P   ,�Ͻ��Ͻ!�Ͻ6�Ͻ��Ͻ?�ϽK�Ͻ!�ϽI�Ͻ)�ϽH�Ͻ=�Ͻ<�Ͻ%�Ͻg�Ͻ!�Ͻ>�Ͻ��Ͻ4�Ͻ^�ϽP   P   6�Ͻ��ϽT�Ͻ��Ͻ_�Ͻn�Ͻj�Ͻ��ϽS�Ͻd�Ͻ(�ϽS�Ͻ�Ͻ��Ͻ��Ͻg�Ͻ-�Ͻb�Ͻ��Ͻ �ϽP   P   +�ϽE�ϽP�Ͻ��Ͻ��Ͻy�Ͻ3�Ͻ"�Ͻ��Ͻ[�Ͻ��Ͻ��Ͻ4�Ͻ��Ͻ��Ͻ%�Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   k�Ͻ�Ͻ�Ͻ��ϽD�Ͻt�Ͻ�Ͻ��Ͻ��ϽZ�Ͻ��Ͻ:�ϽQ�Ͻ4�Ͻ�Ͻ<�ϽS�ϽU�ϽQ�Ͻe�ϽP   P   q�Ͻb�Ͻ��Ͻ'�Ͻg�Ͻ��Ͻ�Ͻ��ϽD�ϽL�Ͻ�Ͻ��Ͻ:�Ͻ��ϽS�Ͻ=�Ͻ��Ͻ*�Ͻ��Ͻ�ϽP   P   ��Ͻ�Ͻl�ϽF�ϽS�ϽR�ϽN�ϽB�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ(�ϽH�ϽJ�Ͻ��ϽX�Ͻ2�ϽP   P   A�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�Ͻ/�Ͻt�Ͻ��Ͻ��ϽL�ϽZ�Ͻ[�Ͻd�Ͻ)�Ͻ�ϽB�Ͻ��ϽM�ϽP   P   ��Ͻm�Ͻ\�Ͻ}�Ͻ��Ͻ_�Ͻ@�Ͻ^�Ͻ��Ͻt�Ͻ��ϽD�Ͻ��Ͻ��ϽS�ϽI�Ͻq�Ͻz�Ͻ5�Ͻ�ϽP   P   4�Ͻ��Ͻ��Ͻ[�Ͻ#�Ͻd�Ͻ��Ͻ��Ͻ^�Ͻ/�ϽB�Ͻ��Ͻ��Ͻ"�Ͻ��Ͻ!�Ͻf�ϽG�Ͻ�Ͻ��ϽP   P   `�ϽB�Ͻ �Ͻ9�Ͻ(�Ͻ�Ͻ.�Ͻ��Ͻ@�Ͻ�ϽN�Ͻ�Ͻ�Ͻ3�Ͻj�ϽK�Ͻt�Ͻ�Ͻc�ϽY�ϽP   P   1�Ͻ��Ͻv�ϽR�Ͻ��Ͻ_�Ͻ�Ͻd�Ͻ_�Ͻ�ϽR�Ͻ��Ͻt�Ͻy�Ͻn�Ͻ?�ϽG�Ͻ��Ͻ��Ͻ>�ϽP   P   �Ͻ��Ͻb�Ͻ��ϽY�Ͻ��Ͻ(�Ͻ#�Ͻ��Ͻ�ϽS�Ͻg�ϽD�Ͻ��Ͻ_�Ͻ��Ͻ�Ͻ:�Ͻ��Ͻ�ϽP   P   T�Ͻd�Ͻ(�Ͻ��Ͻ��ϽR�Ͻ9�Ͻ[�Ͻ}�Ͻ��ϽF�Ͻ'�Ͻ��Ͻ��Ͻ��Ͻ6�Ͻj�ϽW�Ͻ]�Ͻw�ϽP   P   6�Ͻ|�ϽX�Ͻ(�Ͻb�Ͻv�Ͻ �Ͻ��Ͻ\�Ͻ��Ͻl�Ͻ��Ͻ�ϽP�ϽT�Ͻ!�ϽC�Ͻ�Ͻ:�Ͻ�ϽP   P   �ϽB�Ͻ|�Ͻd�Ͻ��Ͻ��ϽB�Ͻ��Ͻm�Ͻ�Ͻ�Ͻb�Ͻ�ϽE�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ(�ϽP   P   ��ϽL�Ͻ8�Ͻ�ϽF�Ͻ[�Ͻ#�Ͻo�Ͻ�Ͻ��Ͻ��Ͻx�Ͻ&�Ͻ��Ͻ8�Ͻ=�Ͻs�Ͻ��Ͻe�ϽV�ϽP   P   V�Ͻ!�ϽB�ϽX�Ͻ��Ͻ^�Ͻ�Ͻ��Ͻi�Ͻ=�ϽR�Ͻl�Ͻ�Ͻi�Ͻ��Ͻ6�Ͻ\�Ͻ��Ͻc�Ͻ�ϽP   P   e�Ͻ��Ͻ\�Ͻd�Ͻ�Ͻ�Ͻ��Ͻ^�Ͻ)�Ͻ��Ͻ\�Ͻ7�Ͻn�Ͻ��Ͻc�ϽU�Ͻ�Ͻ�ϽB�Ͻc�ϽP   P   ��Ͻ��Ͻ-�Ͻ��Ͻ��Ͻ��Ͻ/�Ͻg�Ͻ?�Ͻ�Ͻ��Ͻj�ϽM�Ͻ�Ͻ��Ͻ:�ϽE�ϽY�Ͻ�Ͻ��ϽP   P   s�Ͻ!�Ͻ�Ͻ/�ϽY�ϽM�Ͻ�Ͻo�Ͻ��Ͻ[�Ͻ
�Ͻ��ϽF�Ͻ��ϽI�Ͻ:�Ͻ/�ϽE�Ͻ�Ͻ\�ϽP   P   =�Ͻ��Ͻ=�Ͻ�Ͻ0�Ͻ7�Ͻ2�Ͻ5�ϽC�Ͻc�Ͻ��Ͻ-�ϽK�Ͻc�Ͻ��Ͻ��Ͻ:�Ͻ:�ϽU�Ͻ6�ϽP   P   8�Ͻ��Ͻ6�Ͻ��Ͻ'�Ͻ��Ͻ8�Ͻ��ϽB�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��ϽI�Ͻ��ϽI�Ͻ��Ͻc�Ͻ��ϽP   P   ��Ͻ%�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ-�Ͻo�Ͻ��Ͻ��Ͻ��Ͻ��ϽU�Ͻ-�Ͻ��Ͻc�Ͻ��Ͻ�Ͻ��Ͻi�ϽP   P   &�Ͻ��Ͻ��Ͻ/�ϽJ�Ͻ�Ͻ��Ͻ2�Ͻ�Ͻ-�ϽY�Ͻc�Ͻ)�ϽU�Ͻ�ϽK�ϽF�ϽM�Ͻn�Ͻ�ϽP   P   x�ϽU�Ͻ��ϽG�Ͻ��Ͻ��ϽS�Ͻ��Ͻ`�Ͻ|�Ͻk�Ͻ�Ͻc�Ͻ��Ͻ�Ͻ-�Ͻ��Ͻj�Ͻ7�Ͻl�ϽP   P   ��Ͻ�Ͻ&�Ͻ��Ͻ-�ϽB�Ͻ�Ͻ��Ͻ"�Ͻ>�Ͻ��Ͻk�ϽY�Ͻ��Ͻ�Ͻ��Ͻ
�Ͻ��Ͻ\�ϽR�ϽP   P   ��Ͻ:�Ͻ��Ͻ�Ͻ�Ͻh�Ͻu�Ͻe�Ͻ��Ͻ��Ͻ>�Ͻ|�Ͻ-�Ͻ��Ͻ��Ͻc�Ͻ[�Ͻ�Ͻ��Ͻ=�ϽP   P   �Ͻ@�Ͻ:�Ͻ��Ͻ_�ϽK�ϽX�Ͻi�Ͻf�Ͻ��Ͻ"�Ͻ`�Ͻ�Ͻ��ϽB�ϽC�Ͻ��Ͻ?�Ͻ)�Ͻi�ϽP   P   o�Ͻ<�Ͻ��Ͻ�Ͻ[�Ͻ��Ͻ��Ͻw�Ͻi�Ͻe�Ͻ��Ͻ��Ͻ2�Ͻo�Ͻ��Ͻ5�Ͻo�Ͻg�Ͻ^�Ͻ��ϽP   P   #�Ͻ�Ͻ��ϽC�Ͻ�Ͻo�Ͻ�Ͻ��ϽX�Ͻu�Ͻ�ϽS�Ͻ��Ͻ-�Ͻ8�Ͻ2�Ͻ�Ͻ/�Ͻ��Ͻ�ϽP   P   [�Ͻ��Ͻ�Ͻ.�Ͻ��Ͻ>�Ͻo�Ͻ��ϽK�Ͻh�ϽB�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ7�ϽM�Ͻ��Ͻ�Ͻ^�ϽP   P   F�Ͻ�Ͻ�Ͻ��Ͻ>�Ͻ��Ͻ�Ͻ[�Ͻ_�Ͻ�Ͻ-�Ͻ��ϽJ�Ͻ��Ͻ'�Ͻ0�ϽY�Ͻ��Ͻ�Ͻ��ϽP   P   �Ͻ.�Ͻ>�Ͻ��Ͻ��Ͻ.�ϽC�Ͻ�Ͻ��Ͻ�Ͻ��ϽG�Ͻ/�Ͻ��Ͻ��Ͻ�Ͻ/�Ͻ��Ͻd�ϽX�ϽP   P   8�Ͻ�Ͻ��Ͻ>�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ:�Ͻ��Ͻ&�Ͻ��Ͻ��Ͻ�Ͻ6�Ͻ=�Ͻ�Ͻ-�Ͻ\�ϽB�ϽP   P   L�Ͻs�Ͻ�Ͻ.�Ͻ�Ͻ��Ͻ�Ͻ<�Ͻ@�Ͻ:�Ͻ�ϽU�Ͻ��Ͻ%�Ͻ��Ͻ��Ͻ!�Ͻ��Ͻ��Ͻ!�ϽP   P   ��Ͻ:�Ͻ/�Ͻ��ϽF�Ͻ_�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ:�Ͻ��ϽK�Ͻ2�Ͻ �Ͻ<�Ͻ��Ͻ��Ͻf�Ͻ5�ϽP   P   5�Ͻ��ϽI�Ͻ"�Ͻ��Ͻm�Ͻ	�Ͻ��ϽU�ϽW�Ͻ��Ͻ �Ͻ+�Ͻ*�Ͻ��Ͻ/�ϽR�ϽV�Ͻ%�Ͻ��ϽP   P   f�Ͻ�ϽL�Ͻ�Ͻ$�Ͻ]�Ͻ4�Ͻ9�Ͻ�Ͻw�ϽO�ϽM�Ͻd�Ͻu�Ͻ��Ͻ'�Ͻ^�ϽN�Ͻs�Ͻ%�ϽP   P   ��Ͻ��Ͻ8�Ͻ[�Ͻ��Ͻ`�Ͻ|�Ͻ6�Ͻ�Ͻ��Ͻ}�ϽN�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ�Ͻv�ϽN�ϽV�ϽP   P   ��Ͻa�Ͻ��Ͻ`�Ͻq�ϽR�ϽD�Ͻ(�Ͻ��Ͻ1�Ͻ@�Ͻ[�ϽM�Ͻc�Ͻ��Ͻ�Ͻk�Ͻ�Ͻ^�ϽR�ϽP   P   <�Ͻ��Ͻk�Ͻ,�Ͻ>�Ͻ/�ϽM�Ͻ&�ϽG�Ͻ&�Ͻ��Ͻ��ϽD�Ͻa�ϽT�Ͻ��Ͻ�Ͻ�Ͻ'�Ͻ/�ϽP   P    �Ͻ��ϽC�Ͻ��Ͻ)�Ͻ��Ͻ�Ͻ��Ͻ)�Ͻ��Ͻ`�Ͻy�Ͻ��Ͻ=�Ͻ=�ϽT�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   2�Ͻ��ϽS�Ͻ��Ͻ��ϽB�Ͻ��Ͻ��Ͻc�Ͻ��Ͻ~�Ͻz�Ͻ7�Ͻ��Ͻ=�Ͻa�Ͻc�Ͻ��Ͻu�Ͻ*�ϽP   P   K�Ͻ��Ͻ"�Ͻ�Ͻ>�Ͻ�Ͻ�Ͻ;�Ͻ��Ͻ7�Ͻ7�Ͻ4�Ͻ/�Ͻ7�Ͻ��ϽD�ϽM�Ͻ�Ͻd�Ͻ+�ϽP   P   ��Ͻ��ϽZ�Ͻ.�Ͻ��Ͻp�Ͻb�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ\�Ͻ4�Ͻz�Ͻy�Ͻ��Ͻ[�ϽN�ϽM�Ͻ �ϽP   P   :�ϽP�ϽQ�Ͻ�Ͻ��ϽG�Ͻl�ϽX�Ͻ1�Ͻ[�Ͻ��Ͻ�Ͻ7�Ͻ~�Ͻ`�Ͻ��Ͻ@�Ͻ}�ϽO�Ͻ��ϽP   P   ��ϽL�Ͻx�Ͻ��Ͻ��Ͻ�Ͻ,�Ͻ\�Ͻ��Ͻz�Ͻ[�Ͻ��Ͻ7�Ͻ��Ͻ��Ͻ&�Ͻ1�Ͻ��Ͻw�ϽW�ϽP   P   �Ͻ��ϽR�Ͻ��Ͻ5�Ͻ��Ͻ�Ͻ��Ͻ;�Ͻ��Ͻ1�Ͻ�Ͻ��Ͻc�Ͻ)�ϽG�Ͻ��Ͻ�Ͻ�ϽU�ϽP   P   ��Ͻc�Ͻ,�Ͻ=�Ͻb�Ͻ��ϽK�Ͻ�Ͻ��Ͻ\�ϽX�Ͻ�Ͻ;�Ͻ��Ͻ��Ͻ&�Ͻ(�Ͻ6�Ͻ9�Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻ2�Ͻ�Ͻ*�Ͻ��ϽK�Ͻ�Ͻ,�Ͻl�Ͻb�Ͻ�Ͻ��Ͻ�ϽM�ϽD�Ͻ|�Ͻ4�Ͻ	�ϽP   P   _�Ͻ��ϽX�Ͻ4�Ͻ��Ͻ0�Ͻ*�Ͻ��Ͻ��Ͻ�ϽG�Ͻp�Ͻ�ϽB�Ͻ��Ͻ/�ϽR�Ͻ`�Ͻ]�Ͻm�ϽP   P   F�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ�Ͻb�Ͻ5�Ͻ��Ͻ��Ͻ��Ͻ>�Ͻ��Ͻ)�Ͻ>�Ͻq�Ͻ��Ͻ$�Ͻ��ϽP   P   ��Ͻw�ϽZ�Ͻ��Ͻ��Ͻ4�Ͻ1�Ͻ=�Ͻ��Ͻ��Ͻ�Ͻ.�Ͻ�Ͻ��Ͻ��Ͻ,�Ͻ`�Ͻ[�Ͻ�Ͻ"�ϽP   P   /�Ͻ7�Ͻi�ϽZ�Ͻ�ϽX�Ͻ��Ͻ,�ϽR�Ͻx�ϽQ�ϽZ�Ͻ"�ϽS�ϽC�Ͻk�Ͻ��Ͻ8�ϽL�ϽI�ϽP   P   :�Ͻ�Ͻ7�Ͻw�Ͻ�Ͻ��Ͻ��Ͻc�Ͻ��ϽL�ϽP�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻa�Ͻ��Ͻ�Ͻ��ϽP   P   a�ϽU�Ͻ�Ͻ�Ͻ��Ͻ%�ϽB�Ͻ%�Ͻ��Ͻ��Ͻ �Ͻi�Ͻ��ϽW�Ͻ\�Ͻ�Ͻ��Ͻ�ϽL�Ͻ\�ϽP   P   \�Ͻe�Ͻe�Ͻ+�Ͻ3�Ͻ��Ͻ��ϽW�Ͻ8�Ͻu�Ͻl�Ͻs�Ͻ��Ͻ��Ͻ:�Ͻ��Ͻ��Ͻ�Ͻ
�ϽQ�ϽP   P   L�Ͻ!�ϽB�Ͻ�Ͻ=�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ\�Ͻ	�Ͻ��Ͻ8�Ͻx�ϽO�Ͻ�Ͻf�Ͻ
�ϽP   P   �Ͻ?�ϽN�Ͻ%�Ͻ3�Ͻ3�Ͻ�ϽL�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ(�Ͻ �Ͻ�Ͻ�ϽP   P   ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ"�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ%�Ͻ)�ϽG�Ͻ�Ͻh�Ͻ�Ͻ(�ϽO�Ͻ��ϽP   P   �Ͻ6�Ͻ�Ͻ�ϽD�Ͻ�Ͻ��Ͻ��Ͻ1�Ͻu�Ͻ��ϽT�Ͻ�Ͻ�Ͻ'�Ͻ�Ͻh�Ͻ��Ͻx�Ͻ��ϽP   P   \�Ͻ�Ͻx�Ͻ$�Ͻt�Ͻ�ϽE�Ͻ;�Ͻ��Ͻ��Ͻ �Ͻ5�Ͻp�Ͻ��Ͻ��Ͻ'�Ͻ�Ͻ��Ͻ8�Ͻ:�ϽP   P   W�Ͻ��ϽE�ϽZ�Ͻd�Ͻ0�Ͻ��ϽV�Ͻ$�Ͻ(�Ͻ��Ͻ=�Ͻ�Ͻ.�Ͻ��Ͻ�ϽG�Ͻ��Ͻ��Ͻ��ϽP   P   ��ϽO�Ͻ�Ͻ��Ͻe�Ͻ��Ͻ��Ͻi�Ͻ��ϽY�Ͻ��Ͻ�ϽE�Ͻ�Ͻp�Ͻ�Ͻ)�Ͻ�Ͻ	�Ͻ��ϽP   P   i�Ͻk�Ͻ�Ͻ�Ͻ&�Ͻ �Ͻ3�Ͻ��Ͻ��Ͻ��Ͻk�Ͻi�Ͻ�Ͻ=�Ͻ5�ϽT�Ͻ%�Ͻ�Ͻ\�Ͻs�ϽP   P    �ϽT�Ͻ6�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ.�Ͻ8�Ͻ3�Ͻ�Ͻk�Ͻ��Ͻ��Ͻ �Ͻ��Ͻ��Ͻ��Ͻ��Ͻl�ϽP   P   ��Ͻ-�Ͻ�Ͻ��Ͻ�Ͻ �ϽS�Ͻ��Ͻ��Ͻ�Ͻ3�Ͻ��ϽY�Ͻ(�Ͻ��Ͻu�Ͻ��Ͻ��Ͻ��Ͻu�ϽP   P   ��Ͻ��Ͻ5�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ8�Ͻ��Ͻ��Ͻ$�Ͻ��Ͻ1�Ͻ��Ͻ�Ͻ��Ͻ8�ϽP   P   %�Ͻ�Ͻ��Ͻ �Ͻ��Ͻ��Ͻ=�Ͻ�Ͻ��Ͻ��Ͻ.�Ͻ��Ͻi�ϽV�Ͻ;�Ͻ��Ͻ�ϽL�Ͻ��ϽW�ϽP   P   B�Ͻ�Ͻ��ϽD�Ͻ �ϽY�Ͻ��Ͻ=�Ͻ��ϽS�Ͻ�Ͻ3�Ͻ��Ͻ��ϽE�Ͻ��Ͻ"�Ͻ�Ͻ�Ͻ��ϽP   P   %�Ͻ	�Ͻ2�Ͻ��Ͻ)�Ͻ��ϽY�Ͻ��Ͻ��Ͻ �Ͻ��Ͻ �Ͻ��Ͻ0�Ͻ�Ͻ�Ͻ��Ͻ3�Ͻ��Ͻ��ϽP   P   ��Ͻ>�Ͻj�Ͻw�Ͻ�Ͻ)�Ͻ �Ͻ��Ͻ��Ͻ�Ͻ�Ͻ&�Ͻe�Ͻd�Ͻt�ϽD�Ͻ��Ͻ3�Ͻ=�Ͻ3�ϽP   P   �Ͻ*�Ͻ0�Ͻ�Ͻw�Ͻ��ϽD�Ͻ �Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��ϽZ�Ͻ$�Ͻ�Ͻ��Ͻ%�Ͻ�Ͻ+�ϽP   P   �ϽN�Ͻ��Ͻ0�Ͻj�Ͻ2�Ͻ��Ͻ��Ͻ5�Ͻ�Ͻ6�Ͻ�Ͻ�ϽE�Ͻx�Ͻ�Ͻ�ϽN�ϽB�Ͻe�ϽP   P   U�Ͻ>�ϽN�Ͻ*�Ͻ>�Ͻ	�Ͻ�Ͻ�Ͻ��Ͻ-�ϽT�Ͻk�ϽO�Ͻ��Ͻ�Ͻ6�Ͻ��Ͻ?�Ͻ!�Ͻe�ϽP   P   )�Ͻ��Ͻ�Ͻ(�Ͻ��Ͻo�ϽQ�Ͻ<�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ=�ϽQ�Ͻo�Ͻ��Ͻ'�Ͻ�Ͻ��ϽP   P   ��Ͻ�Ͻ �Ͻu�Ͻc�Ͻ��Ͻ��Ͻ-�Ͻ;�Ͻ��ϽI�Ͻ�Ͻ�Ͻ�Ͻ^�Ͻ��Ͻv�Ͻ��ϽQ�ϽQ�ϽP   P   �Ͻ �Ͻ�Ͻ;�Ͻ�Ͻ+�Ͻ�Ͻ�Ͻ��Ͻo�ϽC�Ͻ�Ͻ(�Ͻo�Ͻ��Ͻ�Ͻ&�ϽE�Ͻ��ϽQ�ϽP   P   '�Ͻt�Ͻ;�ϽU�ϽM�Ͻf�Ͻt�Ͻ+�Ͻ�Ͻ.�Ͻ��Ͻ\�Ͻ��Ͻy�Ͻ\�Ͻ�Ͻ3�ϽD�ϽE�Ͻ��ϽP   P   ��Ͻa�Ͻ�ϽL�Ͻ��Ͻe�Ͻ!�Ͻ�Ͻ��Ͻ�Ͻg�Ͻ8�ϽV�Ͻ9�ϽD�Ͻ�Ͻ��Ͻ3�Ͻ&�Ͻv�ϽP   P   o�Ͻ��Ͻ)�Ͻe�Ͻd�Ͻ��Ͻ��Ͻ�Ͻ+�Ͻ��Ͻ��Ͻ�Ͻ"�Ͻ��Ͻ(�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��ϽP   P   Q�Ͻ��Ͻ�Ͻs�Ͻ�Ͻ��ϽF�Ͻ*�Ͻ��Ͻ*�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ(�ϽD�Ͻ\�Ͻ��Ͻ^�ϽP   P   =�Ͻ+�Ͻ�Ͻ*�Ͻ�Ͻ�Ͻ)�ϽT�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ9�Ͻy�Ͻo�Ͻ�ϽP   P   ��Ͻ;�Ͻ��Ͻ�Ͻ��Ͻ+�Ͻ��Ͻ�Ͻ��Ͻ��ϽW�Ͻa�Ͻ��Ͻ�Ͻ��Ͻ"�ϽV�Ͻ��Ͻ(�Ͻ�ϽP   P   ��Ͻ��Ͻo�Ͻ,�Ͻ�Ͻ��Ͻ*�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ*�Ͻa�Ͻ�Ͻ�Ͻ�Ͻ8�Ͻ\�Ͻ�Ͻ�ϽP   P   �ϽJ�ϽD�Ͻ��Ͻg�Ͻ��Ͻ��Ͻ��ϽY�Ͻ�Ͻ=�Ͻ�ϽW�Ͻ��Ͻ��Ͻ��Ͻg�Ͻ��ϽC�ϽI�ϽP   P   ��Ͻ�Ͻ�Ͻ^�Ͻ8�Ͻ �Ͻ�Ͻ�Ͻb�Ͻ+�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ*�Ͻ��Ͻ�Ͻ.�Ͻo�Ͻ��ϽP   P   ��Ͻ�Ͻ*�Ͻ��ϽU�Ͻ!�Ͻ��Ͻ�Ͻ��Ͻb�ϽY�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ+�Ͻ��Ͻ�Ͻ��Ͻ;�ϽP   P   <�Ͻ�Ͻo�Ͻz�Ͻ9�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ�ϽT�Ͻ*�Ͻ�Ͻ�Ͻ+�Ͻ�Ͻ-�ϽP   P   Q�Ͻ\�Ͻ��Ͻ\�ϽD�Ͻ&�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ*�Ͻ��Ͻ)�ϽF�Ͻ��Ͻ!�Ͻt�Ͻ�Ͻ��ϽP   P   o�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��Ͻ&�Ͻ��Ͻ!�Ͻ �Ͻ��Ͻ��Ͻ+�Ͻ�Ͻ��Ͻ��Ͻe�Ͻf�Ͻ+�Ͻ��ϽP   P   ��Ͻt�Ͻ$�Ͻ3�Ͻ��Ͻ�ϽD�Ͻ9�ϽU�Ͻ8�Ͻg�Ͻ�Ͻ��Ͻ�Ͻ�Ͻd�Ͻ��ϽM�Ͻ�Ͻc�ϽP   P   (�Ͻ��ϽD�ϽC�Ͻ3�Ͻ�Ͻ\�Ͻz�Ͻ��Ͻ^�Ͻ��Ͻ,�Ͻ�Ͻ*�Ͻs�Ͻe�ϽL�ϽU�Ͻ;�Ͻu�ϽP   P   �ϽP�Ͻ��ϽD�Ͻ$�Ͻ�Ͻ��Ͻo�Ͻ*�Ͻ�ϽD�Ͻo�Ͻ��Ͻ�Ͻ�Ͻ)�Ͻ�Ͻ;�Ͻ�Ͻ �ϽP   P   ��ϽP�ϽP�Ͻ��Ͻt�Ͻ��Ͻ\�Ͻ�Ͻ�Ͻ�ϽJ�Ͻ��Ͻ;�Ͻ+�Ͻ��Ͻ��Ͻa�Ͻt�Ͻ �Ͻ�ϽP   P   X�ϽR�ϽA�Ͻ�Ͻ��Ͻ�ϽR�ϽL�Ͻ��Ͻ]�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ8�Ͻ�Ͻ��Ͻ��Ͻ�ϽK�ϽP   P   K�ϽZ�Ͻ�Ͻ4�Ͻ��Ͻ*�Ͻ	�Ͻ��ϽD�Ͻa�ϽI�Ͻ#�Ͻ��Ͻs�Ͻ�Ͻ��Ͻ1�Ͻ�ϽC�Ͻ2�ϽP   P   �Ͻ[�Ͻ8�ϽC�Ͻ�Ͻ�Ͻl�Ͻ8�Ͻ�Ͻ��Ͻ,�Ͻ��Ͻ+�Ͻ��Ͻ��Ͻ%�Ͻ_�Ͻ$�Ͻ��ϽC�ϽP   P   ��Ͻ �Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�ϽN�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ:�Ͻ��Ͻk�Ͻ
�Ͻ$�Ͻ�ϽP   P   ��Ͻ+�Ͻ3�Ͻ)�Ͻ��Ͻ9�Ͻh�ϽW�Ͻ[�Ͻ�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ �Ͻ�Ͻk�Ͻ_�Ͻ1�ϽP   P   �Ͻ��Ͻ��Ͻ*�Ͻ��Ͻ�Ͻ�Ͻ%�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽL�Ͻ��Ͻ �Ͻ��Ͻ%�Ͻ��ϽP   P   8�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��Ͻ:�Ͻ��Ͻ��Ͻ(�Ͻ�ϽH�Ͻ��Ͻ3�Ͻ��ϽL�Ͻ��Ͻ:�Ͻ��Ͻ�ϽP   P   �ϽN�Ͻ��ϽA�Ͻ�Ͻ�Ͻ1�ϽL�Ͻ\�Ͻ��Ͻ$�Ͻ��Ͻ��Ͻ��Ͻ3�Ͻ��Ͻ��Ͻ�Ͻ��Ͻs�ϽP   P   ��Ͻ.�Ͻ��Ͻ��Ͻ��Ͻ'�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ/�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ+�Ͻ��ϽP   P   ��Ͻj�Ͻ��Ͻ��Ͻ��Ͻj�Ͻ��Ͻ�ϽN�Ͻ��Ͻ)�Ͻ �Ͻ��Ͻ��ϽH�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ#�ϽP   P   �Ͻ`�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ^�Ͻ�Ͻ)�Ͻ/�Ͻ$�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ,�ϽI�ϽP   P   ]�Ͻg�ϽP�Ͻ�Ͻ�ϽI�Ͻ+�Ͻ3�Ͻ�Ͻ^�Ͻ^�Ͻ��Ͻ��Ͻ��Ͻ(�Ͻ��Ͻ�Ͻ�Ͻ��Ͻa�ϽP   P   ��Ͻu�Ͻ��Ͻ�Ͻ�Ͻ�Ͻg�Ͻ�Ͻ;�Ͻ�Ͻ��ϽN�Ͻ��Ͻ\�Ͻ��Ͻ��Ͻ[�Ͻ��Ͻ�ϽD�ϽP   P   L�Ͻ��Ͻ��Ͻ��Ͻ<�Ͻ�Ͻ��Ͻ$�Ͻ�Ͻ3�Ͻ��Ͻ�Ͻ�ϽL�Ͻ��Ͻ%�ϽW�ϽN�Ͻ8�Ͻ��ϽP   P   R�Ͻ0�Ͻ/�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻg�Ͻ+�Ͻ�Ͻ��Ͻ��Ͻ1�Ͻ:�Ͻ�Ͻh�Ͻ�Ͻl�Ͻ	�ϽP   P   �Ͻ��Ͻn�Ͻ��Ͻ]�Ͻ�Ͻ�Ͻ�Ͻ�ϽI�Ͻ��Ͻj�Ͻ'�Ͻ�Ͻ��Ͻ�Ͻ9�Ͻ�Ͻ�Ͻ*�ϽP   P   ��Ͻ��ϽF�Ͻ�Ͻ��Ͻ]�Ͻ�Ͻ<�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽP   P   �Ͻ�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��ϽA�Ͻ�Ͻ*�Ͻ)�Ͻ�ϽC�Ͻ4�ϽP   P   A�Ͻ �Ͻ]�Ͻ�ϽF�Ͻn�Ͻ/�Ͻ��Ͻ��ϽP�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ3�Ͻ��Ͻ8�Ͻ�ϽP   P   R�ϽG�Ͻ �Ͻ�Ͻ��Ͻ��Ͻ0�Ͻ��Ͻu�Ͻg�Ͻ`�Ͻj�Ͻ.�ϽN�Ͻ��Ͻ��Ͻ+�Ͻ �Ͻ[�ϽZ�ϽP   P   ��Ͻ�ϽP�Ͻ|�Ͻ��Ͻ&�Ͻ
�Ͻ�Ͻ5�Ͻ��Ͻ'�Ͻ��Ͻ��Ͻ��Ͻ��ϽI�Ͻ1�Ͻv�Ͻ�Ͻ$�ϽP   P   $�Ͻ��Ͻ	�Ͻ��ϽM�Ͻ��Ͻ��Ͻp�Ͻ��Ͻ��Ͻ<�Ͻ7�Ͻ��ϽO�Ͻ��Ͻ��Ͻ�Ͻc�Ͻ"�Ͻ	�ϽP   P   �Ͻ4�Ͻ6�Ͻ$�Ͻ��ϽU�Ͻ0�ϽA�Ͻ�ϽD�Ͻ:�Ͻa�Ͻ;�Ͻ�Ͻ��ϽF�Ͻ�ϽF�ϽU�Ͻ"�ϽP   P   v�Ͻ�Ͻ�ϽF�ϽK�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻw�Ͻ'�Ͻ�Ͻ�Ͻ��Ͻ��ϽF�Ͻc�ϽP   P   1�Ͻ��Ͻ�Ͻ��Ͻ[�Ͻ)�Ͻ�Ͻ��Ͻ*�Ͻl�Ͻl�Ͻ~�Ͻ �ϽN�Ͻi�Ͻl�Ͻ��Ͻ��Ͻ�Ͻ�ϽP   P   I�ϽV�ϽE�ϽI�Ͻ;�Ͻ�Ͻ��Ͻ.�Ͻ��ϽZ�Ͻ2�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻl�Ͻ�ϽF�Ͻ��ϽP   P   ��Ͻ��Ͻ�Ͻf�Ͻ-�Ͻ6�Ͻ��Ͻ��Ͻ��ϽL�ϽW�Ͻ�Ͻ��Ͻ6�Ͻ��Ͻ�Ͻi�Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ#�Ͻ"�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ&�Ͻ��ϽB�ϽF�Ͻ��Ͻ�Ͻ6�Ͻ��ϽN�Ͻ'�Ͻ�ϽO�ϽP   P   ��Ͻ>�Ͻ�Ͻ��Ͻ��Ͻ1�Ͻ�ϽM�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ&�Ͻ��Ͻ��Ͻ��Ͻ �Ͻw�Ͻ;�Ͻ��ϽP   P   ��ϽC�Ͻa�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ"�Ͻ��ϽF�Ͻb�Ͻ��ϽF�Ͻ�Ͻ��Ͻ~�Ͻ��Ͻa�Ͻ7�ϽP   P   '�Ͻ��Ͻ:�Ͻg�Ͻ+�Ͻr�ϽK�Ͻh�Ͻ"�Ͻ��Ͻ��ϽF�Ͻ�ϽB�ϽW�Ͻ2�Ͻl�Ͻ��Ͻ:�Ͻ<�ϽP   P   ��Ͻ��Ͻ:�Ͻ9�ϽF�Ͻ��Ͻd�Ͻd�Ͻ�ϽI�Ͻ��Ͻ��Ͻ��Ͻ��ϽL�ϽZ�Ͻl�Ͻ�ϽD�Ͻ��ϽP   P   5�Ͻ�ϽP�Ͻ��Ͻ9�Ͻ.�Ͻ��Ͻ"�Ͻ�Ͻ�Ͻ"�Ͻ"�Ͻ��Ͻ&�Ͻ��Ͻ��Ͻ*�Ͻ��Ͻ�Ͻ��ϽP   P   �Ͻ�Ͻ`�Ͻm�ϽM�ϽJ�Ͻ%�Ͻ��Ͻ"�Ͻd�Ͻh�Ͻ��ϽM�Ͻ��Ͻ��Ͻ.�Ͻ��Ͻ��ϽA�Ͻp�ϽP   P   
�Ͻ��Ͻ}�Ͻ��Ͻs�Ͻ@�Ͻ%�Ͻ%�Ͻ��Ͻd�ϽK�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ0�Ͻ��ϽP   P   &�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ@�ϽJ�Ͻ.�Ͻ��Ͻr�Ͻ�Ͻ1�Ͻ�Ͻ6�Ͻ�Ͻ)�Ͻ�ϽU�Ͻ��ϽP   P   ��Ͻ;�ϽG�Ͻ��ϽV�Ͻ��Ͻs�ϽM�Ͻ9�ϽF�Ͻ+�Ͻ�Ͻ��Ͻ�Ͻ-�Ͻ;�Ͻ[�ϽK�Ͻ��ϽM�ϽP   P   |�Ͻ@�Ͻ7�Ͻ_�Ͻ��Ͻ��Ͻ��Ͻm�Ͻ��Ͻ9�Ͻg�Ͻ��Ͻ��Ͻ"�Ͻf�ϽI�Ͻ��ϽF�Ͻ$�Ͻ��ϽP   P   P�Ͻ�Ͻ[�Ͻ7�ϽG�Ͻ�Ͻ}�Ͻ`�ϽP�Ͻ:�Ͻ:�Ͻa�Ͻ�Ͻ#�Ͻ�ϽE�Ͻ�Ͻ�Ͻ6�Ͻ	�ϽP   P   �Ͻ��Ͻ�Ͻ@�Ͻ;�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��ϽC�Ͻ>�Ͻ��Ͻ��ϽV�Ͻ��Ͻ�Ͻ4�Ͻ��ϽP   P   ��Ͻ7�ϽE�Ͻ��ϽS�Ͻ�Ͻ�Ͻx�Ͻ�ϽW�Ͻ��Ͻe�Ͻ��ϽP�Ͻ�Ͻ=�Ͻ&�Ͻ��Ͻ�Ͻ-�ϽP   P   -�Ͻ�Ͻk�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ5�Ͻ��Ͻ�Ͻ �Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽT�ϽP   P   �Ͻ"�Ͻ<�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��Ͻu�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ`�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ:�ϽD�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ(�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ%�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ�ϽP   P   &�Ͻ��Ͻ��Ͻ��Ͻ:�Ͻ�Ͻ�Ͻ��Ͻ(�Ͻ��Ͻ�Ͻ_�Ͻ?�Ͻ;�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��ϽP   P   =�Ͻ@�Ͻ�Ͻ��Ͻ/�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ#�ϽG�Ͻ+�Ͻd�ϽN�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�Ͻ�Ͻb�Ͻ3�Ͻ��ϽT�Ͻ8�Ͻs�Ͻ��ϽN�Ͻ��Ͻ%�Ͻ`�Ͻ��ϽP   P   P�Ͻ��Ͻ>�ϽG�ϽO�Ͻ�Ͻ��ϽN�Ͻ�Ͻ��Ͻ��ϽF�ϽH�ϽW�Ͻs�Ͻd�Ͻ;�Ͻ��Ͻ��Ͻ�ϽP   P   ��ϽJ�Ͻ
�Ͻ�Ͻ��Ͻ$�Ͻ$�Ͻc�Ͻ��ϽB�Ͻ�Ͻ��ϽF�ϽH�Ͻ8�Ͻ+�Ͻ?�Ͻ��Ͻ�Ͻ �ϽP   P   e�Ͻ�Ͻ��Ͻ��Ͻ;�ϽD�Ͻ��Ͻ��Ͻ�Ͻ[�Ͻ�Ͻ��Ͻ��ϽF�ϽT�ϽG�Ͻ_�Ͻ��Ͻ��Ͻ�ϽP   P   ��Ͻ1�Ͻ=�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ9�ϽI�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ#�Ͻ�Ͻ��Ͻ�Ͻ��ϽP   P   W�ϽJ�Ͻ�ϽJ�Ͻ��Ͻ�Ͻ��Ͻ��ϽD�Ͻ��ϽI�Ͻ[�ϽB�Ͻ��Ͻ3�Ͻ��Ͻ��Ͻ(�Ͻ��Ͻ5�ϽP   P   �Ͻ��ϽO�Ͻ,�Ͻ'�Ͻ+�Ͻ��Ͻ5�Ͻ�ϽD�Ͻ9�Ͻ�Ͻ��Ͻ�Ͻb�Ͻ��Ͻ(�Ͻ�Ͻu�Ͻ��ϽP   P   x�ϽI�Ͻ��Ͻ��Ͻ��ϽE�Ͻ��Ͻ�Ͻ5�Ͻ��Ͻ��Ͻ��Ͻc�ϽN�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   �Ͻ�ϽC�Ͻ��Ͻ)�Ͻ��Ͻ,�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ$�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��ϽP   P   �Ͻ�Ͻ6�Ͻ�Ͻ�Ͻ��Ͻ��ϽE�Ͻ+�Ͻ�Ͻ��ϽD�Ͻ$�Ͻ�Ͻ�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ��ϽP   P   S�Ͻ=�Ͻ��Ͻ&�Ͻ�Ͻ�Ͻ)�Ͻ��Ͻ'�Ͻ��Ͻ��Ͻ;�Ͻ��ϽO�Ͻ��Ͻ/�Ͻ:�Ͻ�Ͻ��Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻ;�Ͻ&�Ͻ�Ͻ��Ͻ��Ͻ,�ϽJ�Ͻ��Ͻ��Ͻ�ϽG�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽP   P   E�ϽD�Ͻ$�Ͻ��Ͻ��Ͻ6�ϽC�Ͻ��ϽO�Ͻ�Ͻ=�Ͻ��Ͻ
�Ͻ>�Ͻ��Ͻ�Ͻ��ϽD�Ͻ<�Ͻk�ϽP   P   7�Ͻ��ϽD�Ͻ��Ͻ=�Ͻ�Ͻ�ϽI�Ͻ��ϽJ�Ͻ1�Ͻ�ϽJ�Ͻ��Ͻ��Ͻ@�Ͻ��Ͻ:�Ͻ"�Ͻ�ϽP   P   Q�Ͻ��Ͻ�Ͻ �Ͻ��Ͻ�Ͻ�Ͻ�ϽA�ϽG�Ͻm�Ͻ�Ͻa�Ͻ
�Ͻ6�Ͻ�Ͻ��Ͻ+�Ͻ�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻe�ϽX�Ͻu�Ͻr�Ͻ�Ͻ��Ͻ8�Ͻ��Ͻ��ϽC�Ͻ��Ͻ�ϽW�Ͻf�Ͻ:�ϽR�Ͻ�ϽP   P   �Ͻ��Ͻ�ϽU�Ͻ�Ͻ��Ͻ,�Ͻ(�Ͻ��Ͻ��ϽA�Ͻ��Ͻ0�Ͻ��Ͻ��ϽM�Ͻ9�Ͻ��Ͻ.�ϽR�ϽP   P   +�ϽL�Ͻ2�Ͻ.�Ͻ@�Ͻ�Ͻ��Ͻ��Ͻ_�Ͻ��Ͻ�ϽX�ϽQ�Ͻ/�Ͻ�Ͻ)�Ͻ��Ͻ��Ͻ��Ͻ:�ϽP   P   ��Ͻ��Ͻv�Ͻ�Ͻ��ϽY�Ͻ4�Ͻ��Ͻ�Ͻ<�Ͻ(�Ͻ��Ͻ��Ͻ��Ͻ��ϽU�Ͻ0�Ͻ��Ͻ9�Ͻf�ϽP   P   �Ͻ�Ͻv�Ͻg�Ͻ�Ͻ�ϽE�ϽQ�ϽJ�Ͻq�Ͻ'�Ͻ��Ͻ5�Ͻ:�Ͻ��Ͻ4�ϽU�Ͻ)�ϽM�ϽW�ϽP   P   6�Ͻ/�Ͻ7�Ͻ��ϽI�Ͻ!�Ͻ@�Ͻ
�Ͻ��Ͻ��Ͻ#�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�ϽP   P   
�Ͻ��Ͻ��Ͻ�Ͻ;�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ5�Ͻ��Ͻ��Ͻ:�Ͻ��Ͻ/�Ͻ��Ͻ��ϽP   P   a�Ͻ��Ͻ�ϽP�ϽG�Ͻ�Ͻ(�Ͻ��Ͻ|�Ͻ�ϽU�ϽG�Ͻ��Ͻ5�Ͻ�Ͻ5�Ͻ��ϽQ�Ͻ0�ϽC�ϽP   P   �Ͻ#�Ͻ\�Ͻ�Ͻ��Ͻ��Ͻ9�Ͻ.�Ͻ0�Ͻ#�Ͻ��Ͻ��ϽG�Ͻ�Ͻ��Ͻ��Ͻ��ϽX�Ͻ��Ͻ��ϽP   P   m�Ͻ
�Ͻ-�Ͻ��Ͻ�Ͻ�Ͻ��Ͻg�Ͻk�Ͻ��Ͻ��Ͻ��ϽU�Ͻ�Ͻ#�Ͻ'�Ͻ(�Ͻ�ϽA�Ͻ��ϽP   P   G�Ͻ��Ͻ��Ͻ�Ͻo�Ͻ�Ͻ*�Ͻd�Ͻ�Ͻ��Ͻ��Ͻ#�Ͻ�Ͻ��Ͻ��Ͻq�Ͻ<�Ͻ��Ͻ��Ͻ8�ϽP   P   A�Ͻ;�Ͻ&�Ͻ+�Ͻ)�Ͻ�Ͻ��Ͻ
�Ͻ'�Ͻ�Ͻk�Ͻ0�Ͻ|�Ͻ��Ͻ��ϽJ�Ͻ�Ͻ_�Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻf�Ͻh�Ͻ\�Ͻ��Ͻ��Ͻ��Ͻ
�Ͻd�Ͻg�Ͻ.�Ͻ��Ͻ��Ͻ
�ϽQ�Ͻ��Ͻ��Ͻ(�Ͻ�ϽP   P   �Ͻ��Ͻ��Ͻ6�Ͻ�Ͻ=�Ͻ��Ͻ��Ͻ��Ͻ*�Ͻ��Ͻ9�Ͻ(�Ͻ��Ͻ@�ϽE�Ͻ4�Ͻ��Ͻ,�Ͻr�ϽP   P   �Ͻ4�Ͻ	�ϽW�Ͻ�Ͻ��Ͻ=�Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ!�Ͻ�ϽY�Ͻ�Ͻ��Ͻu�ϽP   P   ��Ͻ4�Ͻ�Ͻ-�Ͻ �Ͻ�Ͻ�Ͻ\�Ͻ)�Ͻo�Ͻ�Ͻ��ϽG�Ͻ;�ϽI�Ͻ�Ͻ��Ͻ@�Ͻ�ϽX�ϽP   P    �Ͻ �Ͻ`�Ͻ�Ͻ-�ϽW�Ͻ6�Ͻh�Ͻ+�Ͻ�Ͻ��Ͻ�ϽP�Ͻ�Ͻ��Ͻg�Ͻ�Ͻ.�ϽU�Ͻe�ϽP   P   �Ͻ;�Ͻf�Ͻ`�Ͻ�Ͻ	�Ͻ��Ͻf�Ͻ&�Ͻ��Ͻ-�Ͻ\�Ͻ�Ͻ��Ͻ7�Ͻv�Ͻv�Ͻ2�Ͻ�Ͻ��ϽP   P   ��Ͻ��Ͻ;�Ͻ �Ͻ4�Ͻ4�Ͻ��Ͻ��Ͻ;�Ͻ��Ͻ
�Ͻ#�Ͻ��Ͻ��Ͻ/�Ͻ�Ͻ��ϽL�Ͻ��Ͻ��ϽP   P   ��Ͻ?�Ͻ�Ͻ4�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ6�Ͻ��Ͻ��Ͻ�Ͻ0�Ͻ��Ͻb�ϽF�Ͻ
�Ͻ1�ϽP   P   1�Ͻs�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ@�Ͻ��Ͻ�Ͻ>�ϽV�Ͻ2�Ͻ`�Ͻ(�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   
�Ͻ<�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ �Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽT�Ͻ��Ͻ:�Ͻ+�ϽD�Ͻ��ϽP   P   F�Ͻ��Ͻ��Ͻf�Ͻ��ϽX�ϽZ�Ͻ>�Ͻ�Ͻ1�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ<�Ͻ��Ͻ�Ͻ9�Ͻ+�Ͻ��ϽP   P   b�Ͻ2�Ͻ��Ͻ5�Ͻ#�Ͻ��Ͻ#�Ͻ �Ͻ��Ͻ��Ͻ>�Ͻ
�Ͻ �Ͻ+�Ͻ�Ͻ��Ͻ!�Ͻ�Ͻ:�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ)�Ͻ��Ͻ�Ͻ:�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   0�ϽC�ϽJ�Ͻ��Ͻ/�Ͻ�Ͻ-�Ͻ'�Ͻ8�Ͻ�Ͻ>�Ͻ��ϽV�Ͻ#�Ͻv�Ͻ�Ͻ�Ͻ<�ϽT�Ͻ(�ϽP   P   �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻl�Ͻ6�Ͻq�Ͻ0�Ͻ�Ͻ6�Ͻ#�Ͻ��Ͻ+�Ͻ��Ͻ�Ͻ`�ϽP   P   ��Ͻ�Ͻf�Ͻ��Ͻ�Ͻ��Ͻj�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ	�Ͻ�ϽV�Ͻ)�Ͻ �Ͻ��Ͻ��Ͻ2�ϽP   P   ��Ͻ��ϽQ�Ͻ��Ͻ�Ͻ�ϽA�Ͻ)�Ͻ��Ͻ��Ͻ>�Ͻ��Ͻ��Ͻ0�Ͻ��Ͻ�Ͻ
�Ͻ��Ͻ��ϽV�ϽP   P   6�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��ϽH�Ͻ��Ͻ>�Ͻ��Ͻq�Ͻ>�Ͻ�Ͻ>�Ͻ��Ͻ��Ͻ>�ϽP   P   ��ϽQ�Ͻ��Ͻ��Ͻ3�Ͻ��Ͻ'�Ͻ�Ͻ��Ͻ��ϽH�Ͻ��Ͻ��Ͻ6�Ͻ�Ͻ��Ͻ��Ͻ1�Ͻ��Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻl�Ͻ8�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��ϽP   P   ��Ͻ8�Ͻe�Ͻ��Ͻ)�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ)�Ͻ�Ͻ�Ͻ'�Ͻ�Ͻ �Ͻ>�Ͻ��Ͻ@�ϽP   P   ��Ͻ-�Ͻ��Ͻ7�Ͻ��ϽR�ϽO�Ͻ�Ͻ��Ͻ'�Ͻ�ϽA�Ͻj�Ͻ��Ͻ-�Ͻ��Ͻ#�ϽZ�Ͻ �Ͻ��ϽP   P   ��ϽA�Ͻ�Ͻ �Ͻ8�Ͻ��ϽR�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��ϽX�Ͻ�Ͻ��ϽP   P   ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ8�Ͻ��Ͻ)�Ͻ��Ͻ3�Ͻ�Ͻ�Ͻ�Ͻ��Ͻ/�Ͻ��Ͻ#�Ͻ��Ͻ��Ͻ��ϽP   P   4�Ͻv�Ͻ��Ͻ�Ͻ��Ͻ �Ͻ7�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ5�Ͻf�Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻb�Ͻ��Ͻ��Ͻ�Ͻ��Ͻe�Ͻ��Ͻ��Ͻ��ϽQ�Ͻf�Ͻ��ϽJ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ?�Ͻv�Ͻ��Ͻv�Ͻ�ϽA�Ͻ-�Ͻ8�Ͻ��ϽQ�Ͻ��Ͻ��Ͻ�Ͻ��ϽC�Ͻ��Ͻ2�Ͻ��Ͻ<�Ͻs�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ�ϽT�Ͻ��Ͻ��Ͻ��ϽF�Ͻ��Ͻ
�Ͻ�Ͻ��Ͻ5�Ͻ<�Ͻ_�Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ�ϽF�Ͻ1�Ͻ��Ͻ(�Ͻ
�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ?�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ%�ϽH�ϽP   P   �Ͻ�Ͻ��Ͻ9�Ͻ0�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻ$�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ%�ϽP   P   ��Ͻ3�ϽI�Ͻ��Ͻ��Ͻ��Ͻ�ϽP�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ0�Ͻ��Ͻ��Ͻ��ϽP   P   _�Ͻ��Ͻb�Ͻ �Ͻ�Ͻ�Ͻ��Ͻ4�Ͻ6�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻa�Ͻ0�Ͻ�Ͻ�ϽP   P   <�Ͻ��Ͻ&�Ͻ�Ͻ��ϽT�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ8�Ͻ1�Ͻ��Ͻ��Ͻ�ϽT�Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   5�Ͻ��Ͻ%�ϽK�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ7�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ'�Ͻ�Ͻ.�Ͻa�Ͻ �ϽQ�Ͻ��Ͻ��ϽM�Ͻ��Ͻ��Ͻ��Ͻ.�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ$�Ͻ��ϽP   P   �Ͻ0�Ͻ��Ͻ�Ͻ=�Ͻ��Ͻ��Ͻ6�Ͻ��Ͻ�Ͻ��Ͻ�Ͻr�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�ϽP   P   
�ϽM�Ͻ��Ͻ��Ͻ=�Ͻ0�Ͻ��Ͻ��Ͻj�Ͻ�Ͻ3�Ͻ��Ͻ�Ͻ��Ͻ�Ͻ1�Ͻ��Ͻ��Ͻ��Ͻ?�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻd�Ͻi�ϽF�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ3�Ͻ��Ͻ��Ͻ��Ͻ8�Ͻ��Ͻ��Ͻ�Ͻ�ϽP   P   F�Ͻ��Ͻ��ϽN�Ͻ�Ͻ��Ͻ��Ͻ��ϽW�Ͻ��Ͻ��Ͻ�Ͻ�ϽM�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻ�ϽP   P   ��Ͻ>�Ͻ�Ͻ^�Ͻ�Ͻ��Ͻ
�Ͻ��Ͻ!�ϽW�Ͻ��Ͻj�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ6�Ͻ�Ͻ��Ͻ��ϽP   P   ��ϽZ�Ͻ��Ͻ��Ͻ��Ͻ��ϽS�Ͻ,�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ6�Ͻ��Ͻ��Ͻ��Ͻ4�ϽP�Ͻ��Ͻ��ϽP   P   ��ϽS�Ͻ��Ͻ��ϽS�Ͻ��Ͻ��ϽS�Ͻ
�Ͻ��ϽF�Ͻ��Ͻ��ϽQ�Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ
�ϽP   P   T�Ͻ��Ͻ�Ͻ �ϽW�ϽC�Ͻ��Ͻ��Ͻ��Ͻ��Ͻi�Ͻ0�Ͻ��Ͻ �Ͻ��ϽT�Ͻ�Ͻ��Ͻ��Ͻ(�ϽP   P   �Ͻ��Ͻ��ϽZ�Ͻ��ϽW�ϽS�Ͻ��Ͻ�Ͻ�Ͻd�Ͻ=�Ͻ=�Ͻa�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ0�Ͻ��ϽP   P   ��Ͻ$�Ͻ&�Ͻb�ϽZ�Ͻ �Ͻ��Ͻ��Ͻ^�ϽN�Ͻ��Ͻ��Ͻ�Ͻ.�ϽK�Ͻ�Ͻ �Ͻ��Ͻ9�Ͻ1�ϽP   P   ��Ͻ=�Ͻ?�Ͻ&�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ%�Ͻ&�Ͻb�ϽI�Ͻ��ϽF�ϽP   P   ��Ͻ�Ͻ=�Ͻ$�Ͻ��Ͻ��ϽS�ϽZ�Ͻ>�Ͻ��Ͻ��ϽM�Ͻ0�Ͻ'�Ͻ��Ͻ��Ͻ��Ͻ3�Ͻ�Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��Ͻ&�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ-�Ͻ�Ͻ�ϽQ�Ͻ��Ͻ��Ͻh�Ͻ��Ͻ��Ͻ��ϽI�Ͻ)�Ͻ�Ͻ�Ͻ�Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�Ͻ_�Ͻ �Ͻ��Ͻ`�Ͻ�Ͻe�Ͻ��Ͻ�ϽH�Ͻ�Ͻ �Ͻ��Ͻ�ϽP   P   �Ͻ��Ͻ0�Ͻ��Ͻ2�Ͻ��Ͻ��Ͻ��Ͻ��ϽI�Ͻ�Ͻ�Ͻ��Ͻ �Ͻ�Ͻ�Ͻ��Ͻ��Ͻ �Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ8�Ͻ�Ͻ��Ͻ��ϽI�Ͻ.�Ͻ�Ͻ��Ͻ �Ͻb�Ͻ3�Ͻ��Ͻ��Ͻ�Ͻ�ϽP   P   ��Ͻ%�Ͻ$�Ͻ �ϽT�Ͻ��Ͻ.�ϽS�Ͻ��Ͻ=�Ͻ��Ͻ7�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ3�Ͻ�ϽH�Ͻ)�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻo�Ͻ��ϽL�Ͻ'�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��Ͻb�Ͻ�Ͻ�ϽI�ϽP   P   �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ,�Ͻ��Ͻ1�Ͻ�Ͻ��Ͻ �Ͻ �Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻ��Ͻ<�Ͻ��ϽU�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ%�Ͻ)�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻe�Ͻ��ϽP   P   &�Ͻ�Ͻ��ϽP�Ͻq�Ͻw�ϽR�Ͻ�Ͻ!�Ͻ�Ͻ��Ͻ��Ͻ)�Ͻ,�Ͻ�Ͻ7�Ͻ�Ͻ�Ͻ�Ͻ��ϽP   P   ��Ͻ��ϽX�Ͻ]�Ͻ��Ͻ��Ͻ��Ͻs�Ͻ�Ͻ�Ͻ��Ͻ��Ͻ%�Ͻ�Ͻ'�Ͻ��Ͻ.�Ͻ�Ͻ`�Ͻh�ϽP   P   �Ͻ �Ͻ��Ͻ��Ͻ��ϽH�Ͻ0�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�Ͻ��ϽL�Ͻ=�ϽI�ϽI�Ͻ��Ͻ��ϽP   P   �Ͻ��Ͻ[�Ͻ��Ͻ�Ͻ*�Ͻ��Ͻ/�Ͻ��Ͻ��Ͻ�Ͻ!�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ �Ͻ��ϽP   P   �Ͻ��Ͻ�Ͻ_�Ͻ��Ͻ2�Ͻ��Ͻ��Ͻ/�Ͻ��Ͻs�Ͻ�Ͻ��Ͻ�Ͻo�ϽS�Ͻ��Ͻ��Ͻ_�ϽQ�ϽP   P   ��Ͻ��Ͻ�Ͻ �Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ0�Ͻ��ϽR�Ͻ��Ͻ��Ͻ��Ͻ.�Ͻ�Ͻ��Ͻ�Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻc�Ͻ`�Ͻ��Ͻ�Ͻ2�Ͻ*�ϽH�Ͻ��Ͻw�ϽU�Ͻ��Ͻ��Ͻ��Ͻ8�Ͻ��Ͻ�Ͻ�ϽP   P   ��Ͻ&�Ͻ�Ͻ��Ͻ��Ͻ`�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻq�Ͻ��Ͻ��Ͻ��ϽT�Ͻ��Ͻ2�Ͻ��Ͻ-�ϽP   P   �Ͻ��Ͻ�Ͻ�Ͻ��Ͻc�Ͻ �Ͻ_�Ͻ��Ͻ��Ͻ]�ϽP�Ͻ<�Ͻ��Ͻ��Ͻ �Ͻ��Ͻ��Ͻ�Ͻ��ϽP   P   ��Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ�Ͻ�Ͻ[�Ͻ��ϽX�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ$�Ͻ��Ͻ0�Ͻ��Ͻ��ϽP   P   ��Ͻ��Ͻ�Ͻ��Ͻ&�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ �Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ%�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ �Ͻ8�Ͻ2�Ͻ�Ͻ��Ͻ�Ͻ��Ͻ �Ͻ��Ͻ��Ͻ �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ#�Ͻ?�Ͻ�ϽP   P   �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�Ͻ�Ͻ��Ͻ=�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ?�Ͻ(�Ͻ8�Ͻ��Ͻ��Ͻ�Ͻ �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ�Ͻv�Ͻ��ϽP   P   #�Ͻ��Ͻ��Ͻ(�Ͻ��Ͻ��ϽI�ϽW�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻk�Ͻw�Ͻ�Ͻ�ϽP   P   ��Ͻ�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ<�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻk�Ͻ��Ͻ��ϽP   P   ��Ͻ;�Ͻ��Ͻ��Ͻ,�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻy�Ͻ��Ͻ �Ͻ�Ͻ��ϽT�Ͻ��Ͻ�Ͻ��Ͻ��ϽP   P   ��Ͻ9�Ͻ��Ͻ9�Ͻ�Ͻ3�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��ϽP   P   ��Ͻ@�Ͻ��ϽJ�Ͻ�Ͻ��Ͻ8�Ͻ�Ͻ*�Ͻ��Ͻ��Ͻ�Ͻ-�Ͻ�Ͻ�Ͻ�Ͻ�Ͻ��Ͻ�Ͻ=�ϽP   P   ��Ͻ6�Ͻ��Ͻ��Ͻ-�Ͻ��Ͻ��Ͻ!�Ͻ�Ͻ �Ͻ��Ͻ��Ͻ��Ͻ-�Ͻ��Ͻ �Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P    �Ͻ{�Ͻ��Ͻ��ϽX�Ͻj�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�Ͻ��Ͻ��Ͻ�ϽP   P   ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ%�Ͻ��Ͻ��Ͻ��Ͻ)�Ͻ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻy�Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P   ��Ͻ-�Ͻ��Ͻ��Ͻ��Ͻ'�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ)�Ͻ��Ͻ �Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�ϽP   P    �Ͻ}�Ͻ��Ͻ��Ͻ+�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ�Ͻ*�Ͻ��Ͻ��Ͻ<�Ͻ��Ͻ��Ͻ�ϽP   P   ��Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ[�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ!�Ͻ�Ͻ��Ͻ��Ͻ��ϽW�Ͻ��Ͻ��ϽP   P   �Ͻ�Ͻ7�Ͻ��Ͻ��Ͻ��Ͻ>�Ͻ[�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ8�Ͻ��Ͻ��Ͻ��ϽI�Ͻ �Ͻ��ϽP   P   ��Ͻ�Ͻ��Ͻ��Ͻ>�ϽF�Ͻ��Ͻ��Ͻ��Ͻ'�Ͻ%�Ͻj�Ͻ��Ͻ��Ͻ3�Ͻ��Ͻ��Ͻ��Ͻ�Ͻ��ϽP   P   �Ͻ�ϽY�Ͻ�Ͻx�Ͻ>�Ͻ��Ͻ��Ͻ+�Ͻ��Ͻ��ϽX�Ͻ-�Ͻ�Ͻ�Ͻ,�Ͻ��Ͻ��Ͻ��Ͻ��ϽP   P   2�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��ϽJ�Ͻ9�Ͻ��Ͻ�Ͻ(�Ͻ��Ͻ��ϽP   P   8�Ͻ��Ͻ �Ͻ��ϽY�Ͻ��Ͻ7�Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ��Ͻ8�Ͻ��ϽP   P    �Ͻ�Ͻ��Ͻ��Ͻ�Ͻ�Ͻ�Ͻ�Ͻ}�Ͻ-�Ͻ��Ͻ{�Ͻ6�Ͻ@�Ͻ9�Ͻ;�Ͻ�Ͻ��Ͻ(�Ͻ��ϽP   